module REG_CONTROL #( parameter DATA_WIDTH = 16) (
	current_state,
	counter_ifm,
  reg_write_1,
  reg_write_2,
  reg_write_3,
  reg_write_4,
  reg_write_5,
  reg_write_6,
  reg_write_7,
  reg_write_8,
  reg_write_9,
  reg_write_10,
  reg_write_11,
  reg_write_12,
  reg_write_13,
  reg_write_14,
  reg_write_15,
  reg_write_16,
  reg_write_17,
  reg_write_18,
  reg_write_19,
  reg_write_20,
  reg_write_21,
  reg_write_22,
  reg_write_23,
  reg_write_24,
  reg_write_25,
  reg_write_26,
  reg_write_27,
  reg_write_28,
  reg_write_29,
  reg_write_30,
  reg_write_31,
  reg_write_32,
  reg_write_33,
  reg_write_34,
  reg_write_35,
  reg_write_36,
  reg_write_37,
  reg_write_38,
  reg_write_39,
  reg_write_40,
  reg_write_41,
  reg_write_42,
  reg_write_43,
  reg_write_44,
  reg_write_45,
  reg_write_46,
  reg_write_47,
  reg_write_48,
  reg_write_49,
  reg_write_50,
  reg_write_51,
  reg_write_52,
  reg_write_53,
  reg_write_54,
  reg_write_55,
  reg_write_56,
  reg_write_57,
  reg_write_58,
  reg_write_59,
  reg_write_60,
  reg_write_61,
  reg_write_62,
  reg_write_63,
  reg_write_64,
  reg_write_65,
  reg_write_66,
  reg_write_67,
  reg_write_68,
  reg_write_69,
  reg_write_70,
  reg_write_71,
  reg_write_72,
  reg_write_73,
  reg_write_74,
  reg_write_75,
  reg_write_76,
  reg_write_77,
  reg_write_78,
  reg_write_79,
  reg_write_80,
  reg_write_81,
  reg_write_82,
  reg_write_83,
  reg_write_84,
  reg_write_85,
  reg_write_86,
  reg_write_87,
  reg_write_88,
  reg_write_89,
  reg_write_90,
  reg_write_91,
  reg_write_92,
  reg_write_93,
  reg_write_94,
  reg_write_95,
  reg_write_96,
  reg_write_97,
  reg_write_98,
  reg_write_99,
  reg_write_100,
  reg_write_101,
  reg_write_102,
  reg_write_103,
  reg_write_104,
  reg_write_105,
  reg_write_106,
  reg_write_107,
  reg_write_108,
  reg_write_109,
  reg_write_110,
  reg_write_111,
  reg_write_112,
  reg_write_113,
  reg_write_114,
  reg_write_115,
  reg_write_116,
  reg_write_117,
  reg_write_118,
  reg_write_119,
  reg_write_120,
  reg_write_121,
  reg_write_122,
  reg_write_123,
  reg_write_124,
  reg_write_125,
  reg_write_126,
  reg_write_127,
  reg_write_128,
  reg_write_129,
  reg_write_130,
  reg_write_131,
  reg_write_132,
  reg_write_133,
  reg_write_134,
  reg_write_135,
  reg_write_136,
  reg_write_137,
  reg_write_138,
  reg_write_139,
  reg_write_140,
  reg_write_141,
  reg_write_142,
  reg_write_143,
  reg_write_144,
  reg_write_145,
  reg_write_146,
  reg_write_147,
  reg_write_148,
  reg_write_149,
  reg_write_150,
  reg_write_151,
  reg_write_152,
  reg_write_153,
  reg_write_154,
  reg_write_155,
  reg_write_156,
  reg_write_157,
  reg_write_158,
  reg_write_159,
  reg_write_160,
  reg_write_161,
  reg_write_162,
  reg_write_163,
  reg_write_164,
  reg_write_165,
  reg_write_166,
  reg_write_167,
  reg_write_168,
  reg_write_169,
  reg_write_170,
  reg_write_171,
  reg_write_172,
  reg_write_173,
  reg_write_174,
  reg_write_175,
  reg_write_176,
  reg_write_177,
  reg_write_178,
  reg_write_179,
  reg_write_180,
  reg_write_181,
  reg_write_182,
  reg_write_183,
  reg_write_184,
  reg_write_185,
  reg_write_186,
  reg_write_187,
  reg_write_188,
  reg_write_189,
  reg_write_190,
  reg_write_191,
  reg_write_192,
  reg_write_193,
  reg_write_194,
  reg_write_195,
  reg_write_196,
  reg_write_197,
  reg_write_198,
  reg_write_199,
  reg_write_200,
  reg_write_201,
  reg_write_202,
  reg_write_203,
  reg_write_204,
  reg_write_205,
  reg_write_206,
  reg_write_207,
  reg_write_208,
  reg_write_209,
  reg_write_210,
  reg_write_211,
  reg_write_212,
  reg_write_213,
  reg_write_214,
  reg_write_215,
  reg_write_216,
  reg_write_217,
  reg_write_218,
  reg_write_219,
  reg_write_220,
  reg_write_221,
  reg_write_222,
  reg_write_223,
  reg_write_224,
  reg_write_225,
  reg_write_226,
  reg_write_227,
  reg_write_228,
  reg_write_229,
  reg_write_230,
  reg_write_231,
  reg_write_232,
  reg_write_233,
  reg_write_234,
  reg_write_235,
  reg_write_236,
  reg_write_237,
  reg_write_238,
  reg_write_239,
  reg_write_240,
  reg_write_241,
  reg_write_242,
  reg_write_243,
  reg_write_244,
  reg_write_245,
  reg_write_246,
  reg_write_247,
  reg_write_248,
  reg_write_249,
  reg_write_250,
  reg_write_251,
  reg_write_252,
  reg_write_253,
  reg_write_254,
  reg_write_255,
  reg_write_256,
  reg_write_257,
  reg_write_258,
  reg_write_259,
  reg_write_260,
  reg_write_261,
  reg_write_262,
  reg_write_263,
  reg_write_264,
  reg_write_265,
  reg_write_266,
  reg_write_267,
  reg_write_268,
  reg_write_269,
  reg_write_270,
  reg_write_271,
  reg_write_272,
  reg_write_273,
  reg_write_274,
  reg_write_275,
  reg_write_276,
  reg_write_277,
  reg_write_278,
  reg_write_279,
  reg_write_280,
  reg_write_281,
  reg_write_282,
  reg_write_283,
  reg_write_284,
  reg_write_285,
  reg_write_286,
  reg_write_287,
  reg_write_288,
  reg_write_289,
  reg_write_290,
  reg_write_291,
  reg_write_292,
  reg_write_293,
  reg_write_294,
  reg_write_295,
  reg_write_296,
  reg_write_297,
  reg_write_298,
  reg_write_299,
  reg_write_300,
  reg_write_301,
  reg_write_302,
  reg_write_303,
  reg_write_304,
  reg_write_305,
  reg_write_306,
  reg_write_307,
  reg_write_308,
  reg_write_309,
  reg_write_310,
  reg_write_311,
  reg_write_312,
  reg_write_313,
  reg_write_314,
  reg_write_315,
  reg_write_316,
  reg_write_317,
  reg_write_318,
  reg_write_319,
  reg_write_320,
  reg_write_321,
  reg_write_322,
  reg_write_323,
  reg_write_324,
  reg_write_325,
  reg_write_326,
  reg_write_327,
  reg_write_328,
  reg_write_329,
  reg_write_330,
  reg_write_331,
  reg_write_332,
  reg_write_333,
  reg_write_334,
  reg_write_335,
  reg_write_336,
  reg_write_337,
  reg_write_338,
  reg_write_339,
  reg_write_340,
  reg_write_341,
  reg_write_342,
  reg_write_343,
  reg_write_344,
  reg_write_345,
  reg_write_346,
  reg_write_347,
  reg_write_348,
  reg_write_349,
  reg_write_350,
  reg_write_351,
  reg_write_352,
  reg_write_353,
  reg_write_354,
  reg_write_355,
  reg_write_356,
  reg_write_357,
  reg_write_358,
  reg_write_359,
  reg_write_360,
  reg_write_361,
  reg_write_362,
  reg_write_363,
  reg_write_364,
  reg_write_365,
  reg_write_366,
  reg_write_367,
  reg_write_368,
  reg_write_369,
  reg_write_370,
  reg_write_371,
  reg_write_372,
  reg_write_373,
  reg_write_374,
  reg_write_375,
  reg_write_376,
  reg_write_377,
  reg_write_378,
  reg_write_379,
  reg_write_380,
  reg_write_381,
  reg_write_382,
  reg_write_383,
  reg_write_384,
  reg_write_385,
  reg_write_386,
  reg_write_387,
  reg_write_388,
  reg_write_389,
  reg_write_390,
  reg_write_391,
  reg_write_392,
  reg_write_393,
  reg_write_394,
  reg_write_395,
  reg_write_396,
  reg_write_397,
  reg_write_398,
  reg_write_399,
  reg_write_400,
  reg_write_401,
  reg_write_402,
  reg_write_403,
  reg_write_404,
  reg_write_405,
  reg_write_406,
  reg_write_407,
  reg_write_408,
  reg_write_409,
  reg_write_410,
  reg_write_411,
  reg_write_412,
  reg_write_413,
  reg_write_414,
  reg_write_415,
  reg_write_416,
  reg_write_417,
  reg_write_418,
  reg_write_419,
  reg_write_420,
  reg_write_421,
  reg_write_422,
  reg_write_423,
  reg_write_424,
  reg_write_425,
  reg_write_426,
  reg_write_427,
  reg_write_428,
  reg_write_429,
  reg_write_430,
  reg_write_431,
  reg_write_432,
  reg_write_433,
  reg_write_434,
  reg_write_435,
  reg_write_436,
  reg_write_437,
  reg_write_438,
  reg_write_439,
  reg_write_440,
  reg_write_441,
  reg_write_442,
  reg_write_443,
  reg_write_444,
  reg_write_445,
  reg_write_446,
  reg_write_447,
  reg_write_448,
  reg_write_449,
  reg_write_450,
  reg_write_451,
  reg_write_452,
  reg_write_453,
  reg_write_454,
  reg_write_455,
  reg_write_456,
  reg_write_457,
  reg_write_458,
  reg_write_459,
  reg_write_460,
  reg_write_461,
  reg_write_462,
  reg_write_463,
  reg_write_464,
  reg_write_465,
  reg_write_466,
  reg_write_467,
  reg_write_468,
  reg_write_469,
  reg_write_470,
  reg_write_471,
  reg_write_472,
  reg_write_473,
  reg_write_474,
  reg_write_475,
  reg_write_476,
  reg_write_477,
  reg_write_478,
  reg_write_479,
  reg_write_480,
  reg_write_481,
  reg_write_482,
  reg_write_483,
  reg_write_484,
  reg_write_485,
  reg_write_486,
  reg_write_487,
  reg_write_488,
  reg_write_489,
  reg_write_490,
  reg_write_491,
  reg_write_492,
  reg_write_493,
  reg_write_494,
  reg_write_495,
  reg_write_496,
  reg_write_497,
  reg_write_498,
  reg_write_499,
  reg_write_500,
  reg_write_501,
  reg_write_502,
  reg_write_503,
  reg_write_504,
  reg_write_505,
  reg_write_506,
  reg_write_507,
  reg_write_508,
  reg_write_509,
  reg_write_510,
  reg_write_511,
  reg_write_512,
  reg_write_513,
  reg_write_514,
  reg_write_515,
  reg_write_516,
  reg_write_517,
  reg_write_518,
  reg_write_519,
  reg_write_520,
  reg_write_521,
  reg_write_522,
  reg_write_523,
  reg_write_524,
  reg_write_525,
  reg_write_526,
  reg_write_527,
  reg_write_528,
  reg_write_529,
  reg_write_530,
  reg_write_531,
  reg_write_532,
  reg_write_533,
  reg_write_534,
  reg_write_535,
  reg_write_536,
  reg_write_537,
  reg_write_538,
  reg_write_539,
  reg_write_540,
  reg_write_541,
  reg_write_542,
  reg_write_543,
  reg_write_544,
  reg_write_545,
  reg_write_546,
  reg_write_547,
  reg_write_548,
  reg_write_549,
  reg_write_550,
  reg_write_551,
  reg_write_552,
  reg_write_553,
  reg_write_554,
  reg_write_555,
  reg_write_556,
  reg_write_557,
  reg_write_558,
  reg_write_559,
  reg_write_560,
  reg_write_561,
  reg_write_562,
  reg_write_563,
  reg_write_564,
  reg_write_565,
  reg_write_566,
  reg_write_567,
  reg_write_568,
  reg_write_569,
  reg_write_570,
  reg_write_571,
  reg_write_572,
  reg_write_573,
  reg_write_574,
  reg_write_575,
  reg_write_576,
  reg_write_577,
  reg_write_578,
  reg_write_579,
  reg_write_580,
  reg_write_581,
  reg_write_582,
  reg_write_583,
  reg_write_584,
  reg_write_585,
  reg_write_586,
  reg_write_587,
  reg_write_588,
  reg_write_589,
  reg_write_590,
  reg_write_591,
  reg_write_592,
  reg_write_593,
  reg_write_594,
  reg_write_595,
  reg_write_596,
  reg_write_597,
  reg_write_598,
  reg_write_599,
  reg_write_600,
  reg_write_601,
  reg_write_602,
  reg_write_603,
  reg_write_604,
  reg_write_605,
  reg_write_606,
  reg_write_607,
  reg_write_608,
  reg_write_609,
  reg_write_610,
  reg_write_611,
  reg_write_612,
  reg_write_613,
  reg_write_614,
  reg_write_615,
  reg_write_616,
  reg_write_617,
  reg_write_618,
  reg_write_619,
  reg_write_620,
  reg_write_621,
  reg_write_622,
  reg_write_623,
  reg_write_624,
  reg_write_625,
  reg_write_626,
  reg_write_627,
  reg_write_628,
  reg_write_629,
  reg_write_630,
  reg_write_631,
  reg_write_632,
  reg_write_633,
  reg_write_634,
  reg_write_635,
  reg_write_636,
  reg_write_637,
  reg_write_638,
  reg_write_639,
  reg_write_640,
  reg_write_641,
  reg_write_642,
  reg_write_643,
  reg_write_644,
  reg_write_645,
  reg_write_646,
  reg_write_647,
  reg_write_648,
  reg_write_649,
  reg_write_650,
  reg_write_651,
  reg_write_652,
  reg_write_653,
  reg_write_654,
  reg_write_655,
  reg_write_656,
  reg_write_657,
  reg_write_658,
  reg_write_659,
  reg_write_660,
  reg_write_661,
  reg_write_662,
  reg_write_663,
  reg_write_664,
  reg_write_665,
  reg_write_666,
  reg_write_667,
  reg_write_668,
  reg_write_669,
  reg_write_670,
  reg_write_671,
  reg_write_672,
  reg_write_673,
  reg_write_674,
  reg_write_675,
  reg_write_676,
  reg_write_677,
  reg_write_678,
  reg_write_679,
  reg_write_680,
  reg_write_681,
  reg_write_682,
  reg_write_683,
  reg_write_684,
  reg_write_685,
  reg_write_686,
  reg_write_687,
  reg_write_688,
  reg_write_689,
  reg_write_690,
  reg_write_691,
  reg_write_692,
  reg_write_693,
  reg_write_694,
  reg_write_695,
  reg_write_696,
  reg_write_697,
  reg_write_698,
  reg_write_699,
  reg_write_700,
  reg_write_701,
  reg_write_702,
  reg_write_703,
  reg_write_704,
  reg_write_705,
  reg_write_706,
  reg_write_707,
  reg_write_708,
  reg_write_709,
  reg_write_710,
  reg_write_711,
  reg_write_712,
  reg_write_713,
  reg_write_714,
  reg_write_715,
  reg_write_716,
  reg_write_717,
  reg_write_718,
  reg_write_719,
  reg_write_720,
  reg_write_721,
  reg_write_722,
  reg_write_723,
  reg_write_724,
  reg_write_725,
  reg_write_726,
  reg_write_727,
  reg_write_728,
  reg_write_729,
  reg_write_730,
  reg_write_731,
  reg_write_732,
  reg_write_733,
  reg_write_734,
  reg_write_735,
  reg_write_736,
  reg_write_737,
  reg_write_738,
  reg_write_739,
  reg_write_740,
  reg_write_741,
  reg_write_742,
  reg_write_743,
  reg_write_744,
  reg_write_745,
  reg_write_746,
  reg_write_747,
  reg_write_748,
  reg_write_749,
  reg_write_750,
  reg_write_751,
  reg_write_752,
  reg_write_753,
  reg_write_754,
  reg_write_755,
  reg_write_756,
  reg_write_757,
  reg_write_758,
  reg_write_759,
  reg_write_760,
  reg_write_761,
  reg_write_762,
  reg_write_763,
  reg_write_764,
  reg_write_765,
  reg_write_766,
  reg_write_767,
  reg_write_768,
  reg_write_769,
  reg_write_770,
  reg_write_771,
  reg_write_772,
  reg_write_773,
  reg_write_774,
  reg_write_775,
  reg_write_776,
  reg_write_777,
  reg_write_778,
  reg_write_779,
  reg_write_780,
  reg_write_781,
  reg_write_782,
  reg_write_783,
  reg_write_784,
  reg_write_785,
  reg_write_786,
  reg_write_787,
  reg_write_788,
  reg_write_789,
  reg_write_790,
  reg_write_791,
  reg_write_792,
  reg_write_793,
  reg_write_794,
  reg_write_795,
  reg_write_796,
  reg_write_797,
  reg_write_798,
  reg_write_799,
  reg_write_800,
  reg_write_801,
  reg_write_802,
  reg_write_803,
  reg_write_804,
  reg_write_805,
  reg_write_806,
  reg_write_807,
  reg_write_808,
  reg_write_809,
  reg_write_810,
  reg_write_811,
  reg_write_812,
  reg_write_813,
  reg_write_814,
  reg_write_815,
  reg_write_816,
  reg_write_817,
  reg_write_818,
  reg_write_819,
  reg_write_820,
  reg_write_821,
  reg_write_822,
  reg_write_823,
  reg_write_824,
  reg_write_825,
  reg_write_826,
  reg_write_827,
  reg_write_828,
  reg_write_829,
  reg_write_830,
  reg_write_831,
  reg_write_832,
  reg_write_833,
  reg_write_834,
  reg_write_835,
  reg_write_836,
  reg_write_837,
  reg_write_838,
  reg_write_839,
  reg_write_840,
  reg_write_841,
  reg_write_842,
  reg_write_843,
  reg_write_844,
  reg_write_845,
  reg_write_846,
  reg_write_847,
  reg_write_848,
  reg_write_849,
  reg_write_850,
  reg_write_851,
  reg_write_852,
  reg_write_853,
  reg_write_854,
  reg_write_855,
  reg_write_856,
  reg_write_857,
  reg_write_858,
  reg_write_859,
  reg_write_860,
  reg_write_861,
  reg_write_862,
  reg_write_863,
  reg_write_864,
  reg_write_865,
  reg_write_866,
  reg_write_867,
  reg_write_868,
  reg_write_869,
  reg_write_870,
  reg_write_871,
  reg_write_872,
  reg_write_873,
  reg_write_874,
  reg_write_875,
  reg_write_876,
  reg_write_877,
  reg_write_878,
  reg_write_879,
  reg_write_880,
  reg_write_881,
  reg_write_882,
  reg_write_883,
  reg_write_884,
  reg_write_885,
  reg_write_886,
  reg_write_887,
  reg_write_888,
  reg_write_889,
  reg_write_890,
  reg_write_891,
  reg_write_892,
  reg_write_893,
  reg_write_894,
  reg_write_895,
  reg_write_896,
  reg_write_897,
  reg_write_898,
  reg_write_899,
  reg_write_900,
  reg_write_901,
  reg_write_902,
  reg_write_903,
  reg_write_904,
  reg_write_905,
  reg_write_906,
  reg_write_907,
  reg_write_908,
  reg_write_909,
  reg_write_910,
  reg_write_911,
  reg_write_912,
  reg_write_913,
  reg_write_914,
  reg_write_915,
  reg_write_916,
  reg_write_917,
  reg_write_918,
  reg_write_919,
  reg_write_920,
  reg_write_921,
  reg_write_922,
  reg_write_923,
  reg_write_924,
  reg_write_925,
  reg_write_926,
  reg_write_927,
  reg_write_928,
  reg_write_929,
  reg_write_930,
  reg_write_931,
  reg_write_932,
  reg_write_933,
  reg_write_934,
  reg_write_935,
  reg_write_936,
  reg_write_937,
  reg_write_938,
  reg_write_939,
  reg_write_940,
  reg_write_941,
  reg_write_942,
  reg_write_943,
  reg_write_944,
  reg_write_945,
  reg_write_946,
  reg_write_947,
  reg_write_948,
  reg_write_949,
  reg_write_950,
  reg_write_951,
  reg_write_952,
  reg_write_953,
  reg_write_954,
  reg_write_955,
  reg_write_956,
  reg_write_957,
  reg_write_958,
  reg_write_959,
  reg_write_960,
  reg_write_961,
  reg_write_962,
  reg_write_963,
  reg_write_964,
  reg_write_965,
  reg_write_966,
  reg_write_967,
  reg_write_968,
  reg_write_969,
  reg_write_970,
  reg_write_971,
  reg_write_972,
  reg_write_973,
  reg_write_974,
  reg_write_975,
  reg_write_976,
  reg_write_977,
  reg_write_978,
  reg_write_979,
  reg_write_980,
  reg_write_981,
  reg_write_982,
  reg_write_983,
  reg_write_984,
  reg_write_985,
  reg_write_986,
  reg_write_987,
  reg_write_988,
  reg_write_989,
  reg_write_990,
  reg_write_991,
  reg_write_992,
  reg_write_993,
  reg_write_994,
  reg_write_995,
  reg_write_996,
  reg_write_997,
  reg_write_998,
  reg_write_999,
  reg_write_1000
);

  input [3:0] current_state;
  input [15:0] counter_ifm;
  output reg reg_write_1 ;
  output reg reg_write_2 ;
  output reg reg_write_3 ;
  output reg reg_write_4 ;
  output reg reg_write_5 ;
  output reg reg_write_6 ;
  output reg reg_write_7 ;
  output reg reg_write_8 ;
  output reg reg_write_9 ;
  output reg reg_write_10 ;
  output reg reg_write_11 ;
  output reg reg_write_12 ;
  output reg reg_write_13 ;
  output reg reg_write_14 ;
  output reg reg_write_15 ;
  output reg reg_write_16 ;
  output reg reg_write_17 ;
  output reg reg_write_18 ;
  output reg reg_write_19 ;
  output reg reg_write_20 ;
  output reg reg_write_21 ;
  output reg reg_write_22 ;
  output reg reg_write_23 ;
  output reg reg_write_24 ;
  output reg reg_write_25 ;
  output reg reg_write_26 ;
  output reg reg_write_27 ;
  output reg reg_write_28 ;
  output reg reg_write_29 ;
  output reg reg_write_30 ;
  output reg reg_write_31 ;
  output reg reg_write_32 ;
  output reg reg_write_33 ;
  output reg reg_write_34 ;
  output reg reg_write_35 ;
  output reg reg_write_36 ;
  output reg reg_write_37 ;
  output reg reg_write_38 ;
  output reg reg_write_39 ;
  output reg reg_write_40 ;
  output reg reg_write_41 ;
  output reg reg_write_42 ;
  output reg reg_write_43 ;
  output reg reg_write_44 ;
  output reg reg_write_45 ;
  output reg reg_write_46 ;
  output reg reg_write_47 ;
  output reg reg_write_48 ;
  output reg reg_write_49 ;
  output reg reg_write_50 ;
  output reg reg_write_51 ;
  output reg reg_write_52 ;
  output reg reg_write_53 ;
  output reg reg_write_54 ;
  output reg reg_write_55 ;
  output reg reg_write_56 ;
  output reg reg_write_57 ;
  output reg reg_write_58 ;
  output reg reg_write_59 ;
  output reg reg_write_60 ;
  output reg reg_write_61 ;
  output reg reg_write_62 ;
  output reg reg_write_63 ;
  output reg reg_write_64 ;
  output reg reg_write_65 ;
  output reg reg_write_66 ;
  output reg reg_write_67 ;
  output reg reg_write_68 ;
  output reg reg_write_69 ;
  output reg reg_write_70 ;
  output reg reg_write_71 ;
  output reg reg_write_72 ;
  output reg reg_write_73 ;
  output reg reg_write_74 ;
  output reg reg_write_75 ;
  output reg reg_write_76 ;
  output reg reg_write_77 ;
  output reg reg_write_78 ;
  output reg reg_write_79 ;
  output reg reg_write_80 ;
  output reg reg_write_81 ;
  output reg reg_write_82 ;
  output reg reg_write_83 ;
  output reg reg_write_84 ;
  output reg reg_write_85 ;
  output reg reg_write_86 ;
  output reg reg_write_87 ;
  output reg reg_write_88 ;
  output reg reg_write_89 ;
  output reg reg_write_90 ;
  output reg reg_write_91 ;
  output reg reg_write_92 ;
  output reg reg_write_93 ;
  output reg reg_write_94 ;
  output reg reg_write_95 ;
  output reg reg_write_96 ;
  output reg reg_write_97 ;
  output reg reg_write_98 ;
  output reg reg_write_99 ;
  output reg reg_write_100 ;
  output reg reg_write_101 ;
  output reg reg_write_102 ;
  output reg reg_write_103 ;
  output reg reg_write_104 ;
  output reg reg_write_105 ;
  output reg reg_write_106 ;
  output reg reg_write_107 ;
  output reg reg_write_108 ;
  output reg reg_write_109 ;
  output reg reg_write_110 ;
  output reg reg_write_111 ;
  output reg reg_write_112 ;
  output reg reg_write_113 ;
  output reg reg_write_114 ;
  output reg reg_write_115 ;
  output reg reg_write_116 ;
  output reg reg_write_117 ;
  output reg reg_write_118 ;
  output reg reg_write_119 ;
  output reg reg_write_120 ;
  output reg reg_write_121 ;
  output reg reg_write_122 ;
  output reg reg_write_123 ;
  output reg reg_write_124 ;
  output reg reg_write_125 ;
  output reg reg_write_126 ;
  output reg reg_write_127 ;
  output reg reg_write_128 ;
  output reg reg_write_129 ;
  output reg reg_write_130 ;
  output reg reg_write_131 ;
  output reg reg_write_132 ;
  output reg reg_write_133 ;
  output reg reg_write_134 ;
  output reg reg_write_135 ;
  output reg reg_write_136 ;
  output reg reg_write_137 ;
  output reg reg_write_138 ;
  output reg reg_write_139 ;
  output reg reg_write_140 ;
  output reg reg_write_141 ;
  output reg reg_write_142 ;
  output reg reg_write_143 ;
  output reg reg_write_144 ;
  output reg reg_write_145 ;
  output reg reg_write_146 ;
  output reg reg_write_147 ;
  output reg reg_write_148 ;
  output reg reg_write_149 ;
  output reg reg_write_150 ;
  output reg reg_write_151 ;
  output reg reg_write_152 ;
  output reg reg_write_153 ;
  output reg reg_write_154 ;
  output reg reg_write_155 ;
  output reg reg_write_156 ;
  output reg reg_write_157 ;
  output reg reg_write_158 ;
  output reg reg_write_159 ;
  output reg reg_write_160 ;
  output reg reg_write_161 ;
  output reg reg_write_162 ;
  output reg reg_write_163 ;
  output reg reg_write_164 ;
  output reg reg_write_165 ;
  output reg reg_write_166 ;
  output reg reg_write_167 ;
  output reg reg_write_168 ;
  output reg reg_write_169 ;
  output reg reg_write_170 ;
  output reg reg_write_171 ;
  output reg reg_write_172 ;
  output reg reg_write_173 ;
  output reg reg_write_174 ;
  output reg reg_write_175 ;
  output reg reg_write_176 ;
  output reg reg_write_177 ;
  output reg reg_write_178 ;
  output reg reg_write_179 ;
  output reg reg_write_180 ;
  output reg reg_write_181 ;
  output reg reg_write_182 ;
  output reg reg_write_183 ;
  output reg reg_write_184 ;
  output reg reg_write_185 ;
  output reg reg_write_186 ;
  output reg reg_write_187 ;
  output reg reg_write_188 ;
  output reg reg_write_189 ;
  output reg reg_write_190 ;
  output reg reg_write_191 ;
  output reg reg_write_192 ;
  output reg reg_write_193 ;
  output reg reg_write_194 ;
  output reg reg_write_195 ;
  output reg reg_write_196 ;
  output reg reg_write_197 ;
  output reg reg_write_198 ;
  output reg reg_write_199 ;
  output reg reg_write_200 ;
  output reg reg_write_201 ;
  output reg reg_write_202 ;
  output reg reg_write_203 ;
  output reg reg_write_204 ;
  output reg reg_write_205 ;
  output reg reg_write_206 ;
  output reg reg_write_207 ;
  output reg reg_write_208 ;
  output reg reg_write_209 ;
  output reg reg_write_210 ;
  output reg reg_write_211 ;
  output reg reg_write_212 ;
  output reg reg_write_213 ;
  output reg reg_write_214 ;
  output reg reg_write_215 ;
  output reg reg_write_216 ;
  output reg reg_write_217 ;
  output reg reg_write_218 ;
  output reg reg_write_219 ;
  output reg reg_write_220 ;
  output reg reg_write_221 ;
  output reg reg_write_222 ;
  output reg reg_write_223 ;
  output reg reg_write_224 ;
  output reg reg_write_225 ;
  output reg reg_write_226 ;
  output reg reg_write_227 ;
  output reg reg_write_228 ;
  output reg reg_write_229 ;
  output reg reg_write_230 ;
  output reg reg_write_231 ;
  output reg reg_write_232 ;
  output reg reg_write_233 ;
  output reg reg_write_234 ;
  output reg reg_write_235 ;
  output reg reg_write_236 ;
  output reg reg_write_237 ;
  output reg reg_write_238 ;
  output reg reg_write_239 ;
  output reg reg_write_240 ;
  output reg reg_write_241 ;
  output reg reg_write_242 ;
  output reg reg_write_243 ;
  output reg reg_write_244 ;
  output reg reg_write_245 ;
  output reg reg_write_246 ;
  output reg reg_write_247 ;
  output reg reg_write_248 ;
  output reg reg_write_249 ;
  output reg reg_write_250 ;
  output reg reg_write_251 ;
  output reg reg_write_252 ;
  output reg reg_write_253 ;
  output reg reg_write_254 ;
  output reg reg_write_255 ;
  output reg reg_write_256 ;
  output reg reg_write_257 ;
  output reg reg_write_258 ;
  output reg reg_write_259 ;
  output reg reg_write_260 ;
  output reg reg_write_261 ;
  output reg reg_write_262 ;
  output reg reg_write_263 ;
  output reg reg_write_264 ;
  output reg reg_write_265 ;
  output reg reg_write_266 ;
  output reg reg_write_267 ;
  output reg reg_write_268 ;
  output reg reg_write_269 ;
  output reg reg_write_270 ;
  output reg reg_write_271 ;
  output reg reg_write_272 ;
  output reg reg_write_273 ;
  output reg reg_write_274 ;
  output reg reg_write_275 ;
  output reg reg_write_276 ;
  output reg reg_write_277 ;
  output reg reg_write_278 ;
  output reg reg_write_279 ;
  output reg reg_write_280 ;
  output reg reg_write_281 ;
  output reg reg_write_282 ;
  output reg reg_write_283 ;
  output reg reg_write_284 ;
  output reg reg_write_285 ;
  output reg reg_write_286 ;
  output reg reg_write_287 ;
  output reg reg_write_288 ;
  output reg reg_write_289 ;
  output reg reg_write_290 ;
  output reg reg_write_291 ;
  output reg reg_write_292 ;
  output reg reg_write_293 ;
  output reg reg_write_294 ;
  output reg reg_write_295 ;
  output reg reg_write_296 ;
  output reg reg_write_297 ;
  output reg reg_write_298 ;
  output reg reg_write_299 ;
  output reg reg_write_300 ;
  output reg reg_write_301 ;
  output reg reg_write_302 ;
  output reg reg_write_303 ;
  output reg reg_write_304 ;
  output reg reg_write_305 ;
  output reg reg_write_306 ;
  output reg reg_write_307 ;
  output reg reg_write_308 ;
  output reg reg_write_309 ;
  output reg reg_write_310 ;
  output reg reg_write_311 ;
  output reg reg_write_312 ;
  output reg reg_write_313 ;
  output reg reg_write_314 ;
  output reg reg_write_315 ;
  output reg reg_write_316 ;
  output reg reg_write_317 ;
  output reg reg_write_318 ;
  output reg reg_write_319 ;
  output reg reg_write_320 ;
  output reg reg_write_321 ;
  output reg reg_write_322 ;
  output reg reg_write_323 ;
  output reg reg_write_324 ;
  output reg reg_write_325 ;
  output reg reg_write_326 ;
  output reg reg_write_327 ;
  output reg reg_write_328 ;
  output reg reg_write_329 ;
  output reg reg_write_330 ;
  output reg reg_write_331 ;
  output reg reg_write_332 ;
  output reg reg_write_333 ;
  output reg reg_write_334 ;
  output reg reg_write_335 ;
  output reg reg_write_336 ;
  output reg reg_write_337 ;
  output reg reg_write_338 ;
  output reg reg_write_339 ;
  output reg reg_write_340 ;
  output reg reg_write_341 ;
  output reg reg_write_342 ;
  output reg reg_write_343 ;
  output reg reg_write_344 ;
  output reg reg_write_345 ;
  output reg reg_write_346 ;
  output reg reg_write_347 ;
  output reg reg_write_348 ;
  output reg reg_write_349 ;
  output reg reg_write_350 ;
  output reg reg_write_351 ;
  output reg reg_write_352 ;
  output reg reg_write_353 ;
  output reg reg_write_354 ;
  output reg reg_write_355 ;
  output reg reg_write_356 ;
  output reg reg_write_357 ;
  output reg reg_write_358 ;
  output reg reg_write_359 ;
  output reg reg_write_360 ;
  output reg reg_write_361 ;
  output reg reg_write_362 ;
  output reg reg_write_363 ;
  output reg reg_write_364 ;
  output reg reg_write_365 ;
  output reg reg_write_366 ;
  output reg reg_write_367 ;
  output reg reg_write_368 ;
  output reg reg_write_369 ;
  output reg reg_write_370 ;
  output reg reg_write_371 ;
  output reg reg_write_372 ;
  output reg reg_write_373 ;
  output reg reg_write_374 ;
  output reg reg_write_375 ;
  output reg reg_write_376 ;
  output reg reg_write_377 ;
  output reg reg_write_378 ;
  output reg reg_write_379 ;
  output reg reg_write_380 ;
  output reg reg_write_381 ;
  output reg reg_write_382 ;
  output reg reg_write_383 ;
  output reg reg_write_384 ;
  output reg reg_write_385 ;
  output reg reg_write_386 ;
  output reg reg_write_387 ;
  output reg reg_write_388 ;
  output reg reg_write_389 ;
  output reg reg_write_390 ;
  output reg reg_write_391 ;
  output reg reg_write_392 ;
  output reg reg_write_393 ;
  output reg reg_write_394 ;
  output reg reg_write_395 ;
  output reg reg_write_396 ;
  output reg reg_write_397 ;
  output reg reg_write_398 ;
  output reg reg_write_399 ;
  output reg reg_write_400 ;
  output reg reg_write_401 ;
  output reg reg_write_402 ;
  output reg reg_write_403 ;
  output reg reg_write_404 ;
  output reg reg_write_405 ;
  output reg reg_write_406 ;
  output reg reg_write_407 ;
  output reg reg_write_408 ;
  output reg reg_write_409 ;
  output reg reg_write_410 ;
  output reg reg_write_411 ;
  output reg reg_write_412 ;
  output reg reg_write_413 ;
  output reg reg_write_414 ;
  output reg reg_write_415 ;
  output reg reg_write_416 ;
  output reg reg_write_417 ;
  output reg reg_write_418 ;
  output reg reg_write_419 ;
  output reg reg_write_420 ;
  output reg reg_write_421 ;
  output reg reg_write_422 ;
  output reg reg_write_423 ;
  output reg reg_write_424 ;
  output reg reg_write_425 ;
  output reg reg_write_426 ;
  output reg reg_write_427 ;
  output reg reg_write_428 ;
  output reg reg_write_429 ;
  output reg reg_write_430 ;
  output reg reg_write_431 ;
  output reg reg_write_432 ;
  output reg reg_write_433 ;
  output reg reg_write_434 ;
  output reg reg_write_435 ;
  output reg reg_write_436 ;
  output reg reg_write_437 ;
  output reg reg_write_438 ;
  output reg reg_write_439 ;
  output reg reg_write_440 ;
  output reg reg_write_441 ;
  output reg reg_write_442 ;
  output reg reg_write_443 ;
  output reg reg_write_444 ;
  output reg reg_write_445 ;
  output reg reg_write_446 ;
  output reg reg_write_447 ;
  output reg reg_write_448 ;
  output reg reg_write_449 ;
  output reg reg_write_450 ;
  output reg reg_write_451 ;
  output reg reg_write_452 ;
  output reg reg_write_453 ;
  output reg reg_write_454 ;
  output reg reg_write_455 ;
  output reg reg_write_456 ;
  output reg reg_write_457 ;
  output reg reg_write_458 ;
  output reg reg_write_459 ;
  output reg reg_write_460 ;
  output reg reg_write_461 ;
  output reg reg_write_462 ;
  output reg reg_write_463 ;
  output reg reg_write_464 ;
  output reg reg_write_465 ;
  output reg reg_write_466 ;
  output reg reg_write_467 ;
  output reg reg_write_468 ;
  output reg reg_write_469 ;
  output reg reg_write_470 ;
  output reg reg_write_471 ;
  output reg reg_write_472 ;
  output reg reg_write_473 ;
  output reg reg_write_474 ;
  output reg reg_write_475 ;
  output reg reg_write_476 ;
  output reg reg_write_477 ;
  output reg reg_write_478 ;
  output reg reg_write_479 ;
  output reg reg_write_480 ;
  output reg reg_write_481 ;
  output reg reg_write_482 ;
  output reg reg_write_483 ;
  output reg reg_write_484 ;
  output reg reg_write_485 ;
  output reg reg_write_486 ;
  output reg reg_write_487 ;
  output reg reg_write_488 ;
  output reg reg_write_489 ;
  output reg reg_write_490 ;
  output reg reg_write_491 ;
  output reg reg_write_492 ;
  output reg reg_write_493 ;
  output reg reg_write_494 ;
  output reg reg_write_495 ;
  output reg reg_write_496 ;
  output reg reg_write_497 ;
  output reg reg_write_498 ;
  output reg reg_write_499 ;
  output reg reg_write_500 ;
  output reg reg_write_501 ;
  output reg reg_write_502 ;
  output reg reg_write_503 ;
  output reg reg_write_504 ;
  output reg reg_write_505 ;
  output reg reg_write_506 ;
  output reg reg_write_507 ;
  output reg reg_write_508 ;
  output reg reg_write_509 ;
  output reg reg_write_510 ;
  output reg reg_write_511 ;
  output reg reg_write_512 ;
  output reg reg_write_513 ;
  output reg reg_write_514 ;
  output reg reg_write_515 ;
  output reg reg_write_516 ;
  output reg reg_write_517 ;
  output reg reg_write_518 ;
  output reg reg_write_519 ;
  output reg reg_write_520 ;
  output reg reg_write_521 ;
  output reg reg_write_522 ;
  output reg reg_write_523 ;
  output reg reg_write_524 ;
  output reg reg_write_525 ;
  output reg reg_write_526 ;
  output reg reg_write_527 ;
  output reg reg_write_528 ;
  output reg reg_write_529 ;
  output reg reg_write_530 ;
  output reg reg_write_531 ;
  output reg reg_write_532 ;
  output reg reg_write_533 ;
  output reg reg_write_534 ;
  output reg reg_write_535 ;
  output reg reg_write_536 ;
  output reg reg_write_537 ;
  output reg reg_write_538 ;
  output reg reg_write_539 ;
  output reg reg_write_540 ;
  output reg reg_write_541 ;
  output reg reg_write_542 ;
  output reg reg_write_543 ;
  output reg reg_write_544 ;
  output reg reg_write_545 ;
  output reg reg_write_546 ;
  output reg reg_write_547 ;
  output reg reg_write_548 ;
  output reg reg_write_549 ;
  output reg reg_write_550 ;
  output reg reg_write_551 ;
  output reg reg_write_552 ;
  output reg reg_write_553 ;
  output reg reg_write_554 ;
  output reg reg_write_555 ;
  output reg reg_write_556 ;
  output reg reg_write_557 ;
  output reg reg_write_558 ;
  output reg reg_write_559 ;
  output reg reg_write_560 ;
  output reg reg_write_561 ;
  output reg reg_write_562 ;
  output reg reg_write_563 ;
  output reg reg_write_564 ;
  output reg reg_write_565 ;
  output reg reg_write_566 ;
  output reg reg_write_567 ;
  output reg reg_write_568 ;
  output reg reg_write_569 ;
  output reg reg_write_570 ;
  output reg reg_write_571 ;
  output reg reg_write_572 ;
  output reg reg_write_573 ;
  output reg reg_write_574 ;
  output reg reg_write_575 ;
  output reg reg_write_576 ;
  output reg reg_write_577 ;
  output reg reg_write_578 ;
  output reg reg_write_579 ;
  output reg reg_write_580 ;
  output reg reg_write_581 ;
  output reg reg_write_582 ;
  output reg reg_write_583 ;
  output reg reg_write_584 ;
  output reg reg_write_585 ;
  output reg reg_write_586 ;
  output reg reg_write_587 ;
  output reg reg_write_588 ;
  output reg reg_write_589 ;
  output reg reg_write_590 ;
  output reg reg_write_591 ;
  output reg reg_write_592 ;
  output reg reg_write_593 ;
  output reg reg_write_594 ;
  output reg reg_write_595 ;
  output reg reg_write_596 ;
  output reg reg_write_597 ;
  output reg reg_write_598 ;
  output reg reg_write_599 ;
  output reg reg_write_600 ;
  output reg reg_write_601 ;
  output reg reg_write_602 ;
  output reg reg_write_603 ;
  output reg reg_write_604 ;
  output reg reg_write_605 ;
  output reg reg_write_606 ;
  output reg reg_write_607 ;
  output reg reg_write_608 ;
  output reg reg_write_609 ;
  output reg reg_write_610 ;
  output reg reg_write_611 ;
  output reg reg_write_612 ;
  output reg reg_write_613 ;
  output reg reg_write_614 ;
  output reg reg_write_615 ;
  output reg reg_write_616 ;
  output reg reg_write_617 ;
  output reg reg_write_618 ;
  output reg reg_write_619 ;
  output reg reg_write_620 ;
  output reg reg_write_621 ;
  output reg reg_write_622 ;
  output reg reg_write_623 ;
  output reg reg_write_624 ;
  output reg reg_write_625 ;
  output reg reg_write_626 ;
  output reg reg_write_627 ;
  output reg reg_write_628 ;
  output reg reg_write_629 ;
  output reg reg_write_630 ;
  output reg reg_write_631 ;
  output reg reg_write_632 ;
  output reg reg_write_633 ;
  output reg reg_write_634 ;
  output reg reg_write_635 ;
  output reg reg_write_636 ;
  output reg reg_write_637 ;
  output reg reg_write_638 ;
  output reg reg_write_639 ;
  output reg reg_write_640 ;
  output reg reg_write_641 ;
  output reg reg_write_642 ;
  output reg reg_write_643 ;
  output reg reg_write_644 ;
  output reg reg_write_645 ;
  output reg reg_write_646 ;
  output reg reg_write_647 ;
  output reg reg_write_648 ;
  output reg reg_write_649 ;
  output reg reg_write_650 ;
  output reg reg_write_651 ;
  output reg reg_write_652 ;
  output reg reg_write_653 ;
  output reg reg_write_654 ;
  output reg reg_write_655 ;
  output reg reg_write_656 ;
  output reg reg_write_657 ;
  output reg reg_write_658 ;
  output reg reg_write_659 ;
  output reg reg_write_660 ;
  output reg reg_write_661 ;
  output reg reg_write_662 ;
  output reg reg_write_663 ;
  output reg reg_write_664 ;
  output reg reg_write_665 ;
  output reg reg_write_666 ;
  output reg reg_write_667 ;
  output reg reg_write_668 ;
  output reg reg_write_669 ;
  output reg reg_write_670 ;
  output reg reg_write_671 ;
  output reg reg_write_672 ;
  output reg reg_write_673 ;
  output reg reg_write_674 ;
  output reg reg_write_675 ;
  output reg reg_write_676 ;
  output reg reg_write_677 ;
  output reg reg_write_678 ;
  output reg reg_write_679 ;
  output reg reg_write_680 ;
  output reg reg_write_681 ;
  output reg reg_write_682 ;
  output reg reg_write_683 ;
  output reg reg_write_684 ;
  output reg reg_write_685 ;
  output reg reg_write_686 ;
  output reg reg_write_687 ;
  output reg reg_write_688 ;
  output reg reg_write_689 ;
  output reg reg_write_690 ;
  output reg reg_write_691 ;
  output reg reg_write_692 ;
  output reg reg_write_693 ;
  output reg reg_write_694 ;
  output reg reg_write_695 ;
  output reg reg_write_696 ;
  output reg reg_write_697 ;
  output reg reg_write_698 ;
  output reg reg_write_699 ;
  output reg reg_write_700 ;
  output reg reg_write_701 ;
  output reg reg_write_702 ;
  output reg reg_write_703 ;
  output reg reg_write_704 ;
  output reg reg_write_705 ;
  output reg reg_write_706 ;
  output reg reg_write_707 ;
  output reg reg_write_708 ;
  output reg reg_write_709 ;
  output reg reg_write_710 ;
  output reg reg_write_711 ;
  output reg reg_write_712 ;
  output reg reg_write_713 ;
  output reg reg_write_714 ;
  output reg reg_write_715 ;
  output reg reg_write_716 ;
  output reg reg_write_717 ;
  output reg reg_write_718 ;
  output reg reg_write_719 ;
  output reg reg_write_720 ;
  output reg reg_write_721 ;
  output reg reg_write_722 ;
  output reg reg_write_723 ;
  output reg reg_write_724 ;
  output reg reg_write_725 ;
  output reg reg_write_726 ;
  output reg reg_write_727 ;
  output reg reg_write_728 ;
  output reg reg_write_729 ;
  output reg reg_write_730 ;
  output reg reg_write_731 ;
  output reg reg_write_732 ;
  output reg reg_write_733 ;
  output reg reg_write_734 ;
  output reg reg_write_735 ;
  output reg reg_write_736 ;
  output reg reg_write_737 ;
  output reg reg_write_738 ;
  output reg reg_write_739 ;
  output reg reg_write_740 ;
  output reg reg_write_741 ;
  output reg reg_write_742 ;
  output reg reg_write_743 ;
  output reg reg_write_744 ;
  output reg reg_write_745 ;
  output reg reg_write_746 ;
  output reg reg_write_747 ;
  output reg reg_write_748 ;
  output reg reg_write_749 ;
  output reg reg_write_750 ;
  output reg reg_write_751 ;
  output reg reg_write_752 ;
  output reg reg_write_753 ;
  output reg reg_write_754 ;
  output reg reg_write_755 ;
  output reg reg_write_756 ;
  output reg reg_write_757 ;
  output reg reg_write_758 ;
  output reg reg_write_759 ;
  output reg reg_write_760 ;
  output reg reg_write_761 ;
  output reg reg_write_762 ;
  output reg reg_write_763 ;
  output reg reg_write_764 ;
  output reg reg_write_765 ;
  output reg reg_write_766 ;
  output reg reg_write_767 ;
  output reg reg_write_768 ;
  output reg reg_write_769 ;
  output reg reg_write_770 ;
  output reg reg_write_771 ;
  output reg reg_write_772 ;
  output reg reg_write_773 ;
  output reg reg_write_774 ;
  output reg reg_write_775 ;
  output reg reg_write_776 ;
  output reg reg_write_777 ;
  output reg reg_write_778 ;
  output reg reg_write_779 ;
  output reg reg_write_780 ;
  output reg reg_write_781 ;
  output reg reg_write_782 ;
  output reg reg_write_783 ;
  output reg reg_write_784 ;
  output reg reg_write_785 ;
  output reg reg_write_786 ;
  output reg reg_write_787 ;
  output reg reg_write_788 ;
  output reg reg_write_789 ;
  output reg reg_write_790 ;
  output reg reg_write_791 ;
  output reg reg_write_792 ;
  output reg reg_write_793 ;
  output reg reg_write_794 ;
  output reg reg_write_795 ;
  output reg reg_write_796 ;
  output reg reg_write_797 ;
  output reg reg_write_798 ;
  output reg reg_write_799 ;
  output reg reg_write_800 ;
  output reg reg_write_801 ;
  output reg reg_write_802 ;
  output reg reg_write_803 ;
  output reg reg_write_804 ;
  output reg reg_write_805 ;
  output reg reg_write_806 ;
  output reg reg_write_807 ;
  output reg reg_write_808 ;
  output reg reg_write_809 ;
  output reg reg_write_810 ;
  output reg reg_write_811 ;
  output reg reg_write_812 ;
  output reg reg_write_813 ;
  output reg reg_write_814 ;
  output reg reg_write_815 ;
  output reg reg_write_816 ;
  output reg reg_write_817 ;
  output reg reg_write_818 ;
  output reg reg_write_819 ;
  output reg reg_write_820 ;
  output reg reg_write_821 ;
  output reg reg_write_822 ;
  output reg reg_write_823 ;
  output reg reg_write_824 ;
  output reg reg_write_825 ;
  output reg reg_write_826 ;
  output reg reg_write_827 ;
  output reg reg_write_828 ;
  output reg reg_write_829 ;
  output reg reg_write_830 ;
  output reg reg_write_831 ;
  output reg reg_write_832 ;
  output reg reg_write_833 ;
  output reg reg_write_834 ;
  output reg reg_write_835 ;
  output reg reg_write_836 ;
  output reg reg_write_837 ;
  output reg reg_write_838 ;
  output reg reg_write_839 ;
  output reg reg_write_840 ;
  output reg reg_write_841 ;
  output reg reg_write_842 ;
  output reg reg_write_843 ;
  output reg reg_write_844 ;
  output reg reg_write_845 ;
  output reg reg_write_846 ;
  output reg reg_write_847 ;
  output reg reg_write_848 ;
  output reg reg_write_849 ;
  output reg reg_write_850 ;
  output reg reg_write_851 ;
  output reg reg_write_852 ;
  output reg reg_write_853 ;
  output reg reg_write_854 ;
  output reg reg_write_855 ;
  output reg reg_write_856 ;
  output reg reg_write_857 ;
  output reg reg_write_858 ;
  output reg reg_write_859 ;
  output reg reg_write_860 ;
  output reg reg_write_861 ;
  output reg reg_write_862 ;
  output reg reg_write_863 ;
  output reg reg_write_864 ;
  output reg reg_write_865 ;
  output reg reg_write_866 ;
  output reg reg_write_867 ;
  output reg reg_write_868 ;
  output reg reg_write_869 ;
  output reg reg_write_870 ;
  output reg reg_write_871 ;
  output reg reg_write_872 ;
  output reg reg_write_873 ;
  output reg reg_write_874 ;
  output reg reg_write_875 ;
  output reg reg_write_876 ;
  output reg reg_write_877 ;
  output reg reg_write_878 ;
  output reg reg_write_879 ;
  output reg reg_write_880 ;
  output reg reg_write_881 ;
  output reg reg_write_882 ;
  output reg reg_write_883 ;
  output reg reg_write_884 ;
  output reg reg_write_885 ;
  output reg reg_write_886 ;
  output reg reg_write_887 ;
  output reg reg_write_888 ;
  output reg reg_write_889 ;
  output reg reg_write_890 ;
  output reg reg_write_891 ;
  output reg reg_write_892 ;
  output reg reg_write_893 ;
  output reg reg_write_894 ;
  output reg reg_write_895 ;
  output reg reg_write_896 ;
  output reg reg_write_897 ;
  output reg reg_write_898 ;
  output reg reg_write_899 ;
  output reg reg_write_900 ;
  output reg reg_write_901 ;
  output reg reg_write_902 ;
  output reg reg_write_903 ;
  output reg reg_write_904 ;
  output reg reg_write_905 ;
  output reg reg_write_906 ;
  output reg reg_write_907 ;
  output reg reg_write_908 ;
  output reg reg_write_909 ;
  output reg reg_write_910 ;
  output reg reg_write_911 ;
  output reg reg_write_912 ;
  output reg reg_write_913 ;
  output reg reg_write_914 ;
  output reg reg_write_915 ;
  output reg reg_write_916 ;
  output reg reg_write_917 ;
  output reg reg_write_918 ;
  output reg reg_write_919 ;
  output reg reg_write_920 ;
  output reg reg_write_921 ;
  output reg reg_write_922 ;
  output reg reg_write_923 ;
  output reg reg_write_924 ;
  output reg reg_write_925 ;
  output reg reg_write_926 ;
  output reg reg_write_927 ;
  output reg reg_write_928 ;
  output reg reg_write_929 ;
  output reg reg_write_930 ;
  output reg reg_write_931 ;
  output reg reg_write_932 ;
  output reg reg_write_933 ;
  output reg reg_write_934 ;
  output reg reg_write_935 ;
  output reg reg_write_936 ;
  output reg reg_write_937 ;
  output reg reg_write_938 ;
  output reg reg_write_939 ;
  output reg reg_write_940 ;
  output reg reg_write_941 ;
  output reg reg_write_942 ;
  output reg reg_write_943 ;
  output reg reg_write_944 ;
  output reg reg_write_945 ;
  output reg reg_write_946 ;
  output reg reg_write_947 ;
  output reg reg_write_948 ;
  output reg reg_write_949 ;
  output reg reg_write_950 ;
  output reg reg_write_951 ;
  output reg reg_write_952 ;
  output reg reg_write_953 ;
  output reg reg_write_954 ;
  output reg reg_write_955 ;
  output reg reg_write_956 ;
  output reg reg_write_957 ;
  output reg reg_write_958 ;
  output reg reg_write_959 ;
  output reg reg_write_960 ;
  output reg reg_write_961 ;
  output reg reg_write_962 ;
  output reg reg_write_963 ;
  output reg reg_write_964 ;
  output reg reg_write_965 ;
  output reg reg_write_966 ;
  output reg reg_write_967 ;
  output reg reg_write_968 ;
  output reg reg_write_969 ;
  output reg reg_write_970 ;
  output reg reg_write_971 ;
  output reg reg_write_972 ;
  output reg reg_write_973 ;
  output reg reg_write_974 ;
  output reg reg_write_975 ;
  output reg reg_write_976 ;
  output reg reg_write_977 ;
  output reg reg_write_978 ;
  output reg reg_write_979 ;
  output reg reg_write_980 ;
  output reg reg_write_981 ;
  output reg reg_write_982 ;
  output reg reg_write_983 ;
  output reg reg_write_984 ;
  output reg reg_write_985 ;
  output reg reg_write_986 ;
  output reg reg_write_987 ;
  output reg reg_write_988 ;
  output reg reg_write_989 ;
  output reg reg_write_990 ;
  output reg reg_write_991 ;
  output reg reg_write_992 ;
  output reg reg_write_993 ;
  output reg reg_write_994 ;
  output reg reg_write_995 ;
  output reg reg_write_996 ;
  output reg reg_write_997 ;
  output reg reg_write_998 ;
  output reg reg_write_999 ;
  output reg reg_write_1000 ;

	always @(current_state or counter_ifm) begin
        reg_write_1 = 1'b0 ;
        reg_write_2 = 1'b0 ;
        reg_write_3 = 1'b0 ;
        reg_write_4 = 1'b0 ;
        reg_write_5 = 1'b0 ;
        reg_write_6 = 1'b0 ;
        reg_write_7 = 1'b0 ;
        reg_write_8 = 1'b0 ;
        reg_write_9 = 1'b0 ;
        reg_write_10 = 1'b0 ;
        reg_write_11 = 1'b0 ;
        reg_write_12 = 1'b0 ;
        reg_write_13 = 1'b0 ;
        reg_write_14 = 1'b0 ;
        reg_write_15 = 1'b0 ;
        reg_write_16 = 1'b0 ;
        reg_write_17 = 1'b0 ;
        reg_write_18 = 1'b0 ;
        reg_write_19 = 1'b0 ;
        reg_write_20 = 1'b0 ;
        reg_write_21 = 1'b0 ;
        reg_write_22 = 1'b0 ;
        reg_write_23 = 1'b0 ;
        reg_write_24 = 1'b0 ;
        reg_write_25 = 1'b0 ;
        reg_write_26 = 1'b0 ;
        reg_write_27 = 1'b0 ;
        reg_write_28 = 1'b0 ;
        reg_write_29 = 1'b0 ;
        reg_write_30 = 1'b0 ;
        reg_write_31 = 1'b0 ;
        reg_write_32 = 1'b0 ;
        reg_write_33 = 1'b0 ;
        reg_write_34 = 1'b0 ;
        reg_write_35 = 1'b0 ;
        reg_write_36 = 1'b0 ;
        reg_write_37 = 1'b0 ;
        reg_write_38 = 1'b0 ;
        reg_write_39 = 1'b0 ;
        reg_write_40 = 1'b0 ;
        reg_write_41 = 1'b0 ;
        reg_write_42 = 1'b0 ;
        reg_write_43 = 1'b0 ;
        reg_write_44 = 1'b0 ;
        reg_write_45 = 1'b0 ;
        reg_write_46 = 1'b0 ;
        reg_write_47 = 1'b0 ;
        reg_write_48 = 1'b0 ;
        reg_write_49 = 1'b0 ;
        reg_write_50 = 1'b0 ;
        reg_write_51 = 1'b0 ;
        reg_write_52 = 1'b0 ;
        reg_write_53 = 1'b0 ;
        reg_write_54 = 1'b0 ;
        reg_write_55 = 1'b0 ;
        reg_write_56 = 1'b0 ;
        reg_write_57 = 1'b0 ;
        reg_write_58 = 1'b0 ;
        reg_write_59 = 1'b0 ;
        reg_write_60 = 1'b0 ;
        reg_write_61 = 1'b0 ;
        reg_write_62 = 1'b0 ;
        reg_write_63 = 1'b0 ;
        reg_write_64 = 1'b0 ;
        reg_write_65 = 1'b0 ;
        reg_write_66 = 1'b0 ;
        reg_write_67 = 1'b0 ;
        reg_write_68 = 1'b0 ;
        reg_write_69 = 1'b0 ;
        reg_write_70 = 1'b0 ;
        reg_write_71 = 1'b0 ;
        reg_write_72 = 1'b0 ;
        reg_write_73 = 1'b0 ;
        reg_write_74 = 1'b0 ;
        reg_write_75 = 1'b0 ;
        reg_write_76 = 1'b0 ;
        reg_write_77 = 1'b0 ;
        reg_write_78 = 1'b0 ;
        reg_write_79 = 1'b0 ;
        reg_write_80 = 1'b0 ;
        reg_write_81 = 1'b0 ;
        reg_write_82 = 1'b0 ;
        reg_write_83 = 1'b0 ;
        reg_write_84 = 1'b0 ;
        reg_write_85 = 1'b0 ;
        reg_write_86 = 1'b0 ;
        reg_write_87 = 1'b0 ;
        reg_write_88 = 1'b0 ;
        reg_write_89 = 1'b0 ;
        reg_write_90 = 1'b0 ;
        reg_write_91 = 1'b0 ;
        reg_write_92 = 1'b0 ;
        reg_write_93 = 1'b0 ;
        reg_write_94 = 1'b0 ;
        reg_write_95 = 1'b0 ;
        reg_write_96 = 1'b0 ;
        reg_write_97 = 1'b0 ;
        reg_write_98 = 1'b0 ;
        reg_write_99 = 1'b0 ;
        reg_write_100 = 1'b0 ;
        reg_write_101 = 1'b0 ;
        reg_write_102 = 1'b0 ;
        reg_write_103 = 1'b0 ;
        reg_write_104 = 1'b0 ;
        reg_write_105 = 1'b0 ;
        reg_write_106 = 1'b0 ;
        reg_write_107 = 1'b0 ;
        reg_write_108 = 1'b0 ;
        reg_write_109 = 1'b0 ;
        reg_write_110 = 1'b0 ;
        reg_write_111 = 1'b0 ;
        reg_write_112 = 1'b0 ;
        reg_write_113 = 1'b0 ;
        reg_write_114 = 1'b0 ;
        reg_write_115 = 1'b0 ;
        reg_write_116 = 1'b0 ;
        reg_write_117 = 1'b0 ;
        reg_write_118 = 1'b0 ;
        reg_write_119 = 1'b0 ;
        reg_write_120 = 1'b0 ;
        reg_write_121 = 1'b0 ;
        reg_write_122 = 1'b0 ;
        reg_write_123 = 1'b0 ;
        reg_write_124 = 1'b0 ;
        reg_write_125 = 1'b0 ;
        reg_write_126 = 1'b0 ;
        reg_write_127 = 1'b0 ;
        reg_write_128 = 1'b0 ;
        reg_write_129 = 1'b0 ;
        reg_write_130 = 1'b0 ;
        reg_write_131 = 1'b0 ;
        reg_write_132 = 1'b0 ;
        reg_write_133 = 1'b0 ;
        reg_write_134 = 1'b0 ;
        reg_write_135 = 1'b0 ;
        reg_write_136 = 1'b0 ;
        reg_write_137 = 1'b0 ;
        reg_write_138 = 1'b0 ;
        reg_write_139 = 1'b0 ;
        reg_write_140 = 1'b0 ;
        reg_write_141 = 1'b0 ;
        reg_write_142 = 1'b0 ;
        reg_write_143 = 1'b0 ;
        reg_write_144 = 1'b0 ;
        reg_write_145 = 1'b0 ;
        reg_write_146 = 1'b0 ;
        reg_write_147 = 1'b0 ;
        reg_write_148 = 1'b0 ;
        reg_write_149 = 1'b0 ;
        reg_write_150 = 1'b0 ;
        reg_write_151 = 1'b0 ;
        reg_write_152 = 1'b0 ;
        reg_write_153 = 1'b0 ;
        reg_write_154 = 1'b0 ;
        reg_write_155 = 1'b0 ;
        reg_write_156 = 1'b0 ;
        reg_write_157 = 1'b0 ;
        reg_write_158 = 1'b0 ;
        reg_write_159 = 1'b0 ;
        reg_write_160 = 1'b0 ;
        reg_write_161 = 1'b0 ;
        reg_write_162 = 1'b0 ;
        reg_write_163 = 1'b0 ;
        reg_write_164 = 1'b0 ;
        reg_write_165 = 1'b0 ;
        reg_write_166 = 1'b0 ;
        reg_write_167 = 1'b0 ;
        reg_write_168 = 1'b0 ;
        reg_write_169 = 1'b0 ;
        reg_write_170 = 1'b0 ;
        reg_write_171 = 1'b0 ;
        reg_write_172 = 1'b0 ;
        reg_write_173 = 1'b0 ;
        reg_write_174 = 1'b0 ;
        reg_write_175 = 1'b0 ;
        reg_write_176 = 1'b0 ;
        reg_write_177 = 1'b0 ;
        reg_write_178 = 1'b0 ;
        reg_write_179 = 1'b0 ;
        reg_write_180 = 1'b0 ;
        reg_write_181 = 1'b0 ;
        reg_write_182 = 1'b0 ;
        reg_write_183 = 1'b0 ;
        reg_write_184 = 1'b0 ;
        reg_write_185 = 1'b0 ;
        reg_write_186 = 1'b0 ;
        reg_write_187 = 1'b0 ;
        reg_write_188 = 1'b0 ;
        reg_write_189 = 1'b0 ;
        reg_write_190 = 1'b0 ;
        reg_write_191 = 1'b0 ;
        reg_write_192 = 1'b0 ;
        reg_write_193 = 1'b0 ;
        reg_write_194 = 1'b0 ;
        reg_write_195 = 1'b0 ;
        reg_write_196 = 1'b0 ;
        reg_write_197 = 1'b0 ;
        reg_write_198 = 1'b0 ;
        reg_write_199 = 1'b0 ;
        reg_write_200 = 1'b0 ;
        reg_write_201 = 1'b0 ;
        reg_write_202 = 1'b0 ;
        reg_write_203 = 1'b0 ;
        reg_write_204 = 1'b0 ;
        reg_write_205 = 1'b0 ;
        reg_write_206 = 1'b0 ;
        reg_write_207 = 1'b0 ;
        reg_write_208 = 1'b0 ;
        reg_write_209 = 1'b0 ;
        reg_write_210 = 1'b0 ;
        reg_write_211 = 1'b0 ;
        reg_write_212 = 1'b0 ;
        reg_write_213 = 1'b0 ;
        reg_write_214 = 1'b0 ;
        reg_write_215 = 1'b0 ;
        reg_write_216 = 1'b0 ;
        reg_write_217 = 1'b0 ;
        reg_write_218 = 1'b0 ;
        reg_write_219 = 1'b0 ;
        reg_write_220 = 1'b0 ;
        reg_write_221 = 1'b0 ;
        reg_write_222 = 1'b0 ;
        reg_write_223 = 1'b0 ;
        reg_write_224 = 1'b0 ;
        reg_write_225 = 1'b0 ;
        reg_write_226 = 1'b0 ;
        reg_write_227 = 1'b0 ;
        reg_write_228 = 1'b0 ;
        reg_write_229 = 1'b0 ;
        reg_write_230 = 1'b0 ;
        reg_write_231 = 1'b0 ;
        reg_write_232 = 1'b0 ;
        reg_write_233 = 1'b0 ;
        reg_write_234 = 1'b0 ;
        reg_write_235 = 1'b0 ;
        reg_write_236 = 1'b0 ;
        reg_write_237 = 1'b0 ;
        reg_write_238 = 1'b0 ;
        reg_write_239 = 1'b0 ;
        reg_write_240 = 1'b0 ;
        reg_write_241 = 1'b0 ;
        reg_write_242 = 1'b0 ;
        reg_write_243 = 1'b0 ;
        reg_write_244 = 1'b0 ;
        reg_write_245 = 1'b0 ;
        reg_write_246 = 1'b0 ;
        reg_write_247 = 1'b0 ;
        reg_write_248 = 1'b0 ;
        reg_write_249 = 1'b0 ;
        reg_write_250 = 1'b0 ;
        reg_write_251 = 1'b0 ;
        reg_write_252 = 1'b0 ;
        reg_write_253 = 1'b0 ;
        reg_write_254 = 1'b0 ;
        reg_write_255 = 1'b0 ;
        reg_write_256 = 1'b0 ;
        reg_write_257 = 1'b0 ;
        reg_write_258 = 1'b0 ;
        reg_write_259 = 1'b0 ;
        reg_write_260 = 1'b0 ;
        reg_write_261 = 1'b0 ;
        reg_write_262 = 1'b0 ;
        reg_write_263 = 1'b0 ;
        reg_write_264 = 1'b0 ;
        reg_write_265 = 1'b0 ;
        reg_write_266 = 1'b0 ;
        reg_write_267 = 1'b0 ;
        reg_write_268 = 1'b0 ;
        reg_write_269 = 1'b0 ;
        reg_write_270 = 1'b0 ;
        reg_write_271 = 1'b0 ;
        reg_write_272 = 1'b0 ;
        reg_write_273 = 1'b0 ;
        reg_write_274 = 1'b0 ;
        reg_write_275 = 1'b0 ;
        reg_write_276 = 1'b0 ;
        reg_write_277 = 1'b0 ;
        reg_write_278 = 1'b0 ;
        reg_write_279 = 1'b0 ;
        reg_write_280 = 1'b0 ;
        reg_write_281 = 1'b0 ;
        reg_write_282 = 1'b0 ;
        reg_write_283 = 1'b0 ;
        reg_write_284 = 1'b0 ;
        reg_write_285 = 1'b0 ;
        reg_write_286 = 1'b0 ;
        reg_write_287 = 1'b0 ;
        reg_write_288 = 1'b0 ;
        reg_write_289 = 1'b0 ;
        reg_write_290 = 1'b0 ;
        reg_write_291 = 1'b0 ;
        reg_write_292 = 1'b0 ;
        reg_write_293 = 1'b0 ;
        reg_write_294 = 1'b0 ;
        reg_write_295 = 1'b0 ;
        reg_write_296 = 1'b0 ;
        reg_write_297 = 1'b0 ;
        reg_write_298 = 1'b0 ;
        reg_write_299 = 1'b0 ;
        reg_write_300 = 1'b0 ;
        reg_write_301 = 1'b0 ;
        reg_write_302 = 1'b0 ;
        reg_write_303 = 1'b0 ;
        reg_write_304 = 1'b0 ;
        reg_write_305 = 1'b0 ;
        reg_write_306 = 1'b0 ;
        reg_write_307 = 1'b0 ;
        reg_write_308 = 1'b0 ;
        reg_write_309 = 1'b0 ;
        reg_write_310 = 1'b0 ;
        reg_write_311 = 1'b0 ;
        reg_write_312 = 1'b0 ;
        reg_write_313 = 1'b0 ;
        reg_write_314 = 1'b0 ;
        reg_write_315 = 1'b0 ;
        reg_write_316 = 1'b0 ;
        reg_write_317 = 1'b0 ;
        reg_write_318 = 1'b0 ;
        reg_write_319 = 1'b0 ;
        reg_write_320 = 1'b0 ;
        reg_write_321 = 1'b0 ;
        reg_write_322 = 1'b0 ;
        reg_write_323 = 1'b0 ;
        reg_write_324 = 1'b0 ;
        reg_write_325 = 1'b0 ;
        reg_write_326 = 1'b0 ;
        reg_write_327 = 1'b0 ;
        reg_write_328 = 1'b0 ;
        reg_write_329 = 1'b0 ;
        reg_write_330 = 1'b0 ;
        reg_write_331 = 1'b0 ;
        reg_write_332 = 1'b0 ;
        reg_write_333 = 1'b0 ;
        reg_write_334 = 1'b0 ;
        reg_write_335 = 1'b0 ;
        reg_write_336 = 1'b0 ;
        reg_write_337 = 1'b0 ;
        reg_write_338 = 1'b0 ;
        reg_write_339 = 1'b0 ;
        reg_write_340 = 1'b0 ;
        reg_write_341 = 1'b0 ;
        reg_write_342 = 1'b0 ;
        reg_write_343 = 1'b0 ;
        reg_write_344 = 1'b0 ;
        reg_write_345 = 1'b0 ;
        reg_write_346 = 1'b0 ;
        reg_write_347 = 1'b0 ;
        reg_write_348 = 1'b0 ;
        reg_write_349 = 1'b0 ;
        reg_write_350 = 1'b0 ;
        reg_write_351 = 1'b0 ;
        reg_write_352 = 1'b0 ;
        reg_write_353 = 1'b0 ;
        reg_write_354 = 1'b0 ;
        reg_write_355 = 1'b0 ;
        reg_write_356 = 1'b0 ;
        reg_write_357 = 1'b0 ;
        reg_write_358 = 1'b0 ;
        reg_write_359 = 1'b0 ;
        reg_write_360 = 1'b0 ;
        reg_write_361 = 1'b0 ;
        reg_write_362 = 1'b0 ;
        reg_write_363 = 1'b0 ;
        reg_write_364 = 1'b0 ;
        reg_write_365 = 1'b0 ;
        reg_write_366 = 1'b0 ;
        reg_write_367 = 1'b0 ;
        reg_write_368 = 1'b0 ;
        reg_write_369 = 1'b0 ;
        reg_write_370 = 1'b0 ;
        reg_write_371 = 1'b0 ;
        reg_write_372 = 1'b0 ;
        reg_write_373 = 1'b0 ;
        reg_write_374 = 1'b0 ;
        reg_write_375 = 1'b0 ;
        reg_write_376 = 1'b0 ;
        reg_write_377 = 1'b0 ;
        reg_write_378 = 1'b0 ;
        reg_write_379 = 1'b0 ;
        reg_write_380 = 1'b0 ;
        reg_write_381 = 1'b0 ;
        reg_write_382 = 1'b0 ;
        reg_write_383 = 1'b0 ;
        reg_write_384 = 1'b0 ;
        reg_write_385 = 1'b0 ;
        reg_write_386 = 1'b0 ;
        reg_write_387 = 1'b0 ;
        reg_write_388 = 1'b0 ;
        reg_write_389 = 1'b0 ;
        reg_write_390 = 1'b0 ;
        reg_write_391 = 1'b0 ;
        reg_write_392 = 1'b0 ;
        reg_write_393 = 1'b0 ;
        reg_write_394 = 1'b0 ;
        reg_write_395 = 1'b0 ;
        reg_write_396 = 1'b0 ;
        reg_write_397 = 1'b0 ;
        reg_write_398 = 1'b0 ;
        reg_write_399 = 1'b0 ;
        reg_write_400 = 1'b0 ;
        reg_write_401 = 1'b0 ;
        reg_write_402 = 1'b0 ;
        reg_write_403 = 1'b0 ;
        reg_write_404 = 1'b0 ;
        reg_write_405 = 1'b0 ;
        reg_write_406 = 1'b0 ;
        reg_write_407 = 1'b0 ;
        reg_write_408 = 1'b0 ;
        reg_write_409 = 1'b0 ;
        reg_write_410 = 1'b0 ;
        reg_write_411 = 1'b0 ;
        reg_write_412 = 1'b0 ;
        reg_write_413 = 1'b0 ;
        reg_write_414 = 1'b0 ;
        reg_write_415 = 1'b0 ;
        reg_write_416 = 1'b0 ;
        reg_write_417 = 1'b0 ;
        reg_write_418 = 1'b0 ;
        reg_write_419 = 1'b0 ;
        reg_write_420 = 1'b0 ;
        reg_write_421 = 1'b0 ;
        reg_write_422 = 1'b0 ;
        reg_write_423 = 1'b0 ;
        reg_write_424 = 1'b0 ;
        reg_write_425 = 1'b0 ;
        reg_write_426 = 1'b0 ;
        reg_write_427 = 1'b0 ;
        reg_write_428 = 1'b0 ;
        reg_write_429 = 1'b0 ;
        reg_write_430 = 1'b0 ;
        reg_write_431 = 1'b0 ;
        reg_write_432 = 1'b0 ;
        reg_write_433 = 1'b0 ;
        reg_write_434 = 1'b0 ;
        reg_write_435 = 1'b0 ;
        reg_write_436 = 1'b0 ;
        reg_write_437 = 1'b0 ;
        reg_write_438 = 1'b0 ;
        reg_write_439 = 1'b0 ;
        reg_write_440 = 1'b0 ;
        reg_write_441 = 1'b0 ;
        reg_write_442 = 1'b0 ;
        reg_write_443 = 1'b0 ;
        reg_write_444 = 1'b0 ;
        reg_write_445 = 1'b0 ;
        reg_write_446 = 1'b0 ;
        reg_write_447 = 1'b0 ;
        reg_write_448 = 1'b0 ;
        reg_write_449 = 1'b0 ;
        reg_write_450 = 1'b0 ;
        reg_write_451 = 1'b0 ;
        reg_write_452 = 1'b0 ;
        reg_write_453 = 1'b0 ;
        reg_write_454 = 1'b0 ;
        reg_write_455 = 1'b0 ;
        reg_write_456 = 1'b0 ;
        reg_write_457 = 1'b0 ;
        reg_write_458 = 1'b0 ;
        reg_write_459 = 1'b0 ;
        reg_write_460 = 1'b0 ;
        reg_write_461 = 1'b0 ;
        reg_write_462 = 1'b0 ;
        reg_write_463 = 1'b0 ;
        reg_write_464 = 1'b0 ;
        reg_write_465 = 1'b0 ;
        reg_write_466 = 1'b0 ;
        reg_write_467 = 1'b0 ;
        reg_write_468 = 1'b0 ;
        reg_write_469 = 1'b0 ;
        reg_write_470 = 1'b0 ;
        reg_write_471 = 1'b0 ;
        reg_write_472 = 1'b0 ;
        reg_write_473 = 1'b0 ;
        reg_write_474 = 1'b0 ;
        reg_write_475 = 1'b0 ;
        reg_write_476 = 1'b0 ;
        reg_write_477 = 1'b0 ;
        reg_write_478 = 1'b0 ;
        reg_write_479 = 1'b0 ;
        reg_write_480 = 1'b0 ;
        reg_write_481 = 1'b0 ;
        reg_write_482 = 1'b0 ;
        reg_write_483 = 1'b0 ;
        reg_write_484 = 1'b0 ;
        reg_write_485 = 1'b0 ;
        reg_write_486 = 1'b0 ;
        reg_write_487 = 1'b0 ;
        reg_write_488 = 1'b0 ;
        reg_write_489 = 1'b0 ;
        reg_write_490 = 1'b0 ;
        reg_write_491 = 1'b0 ;
        reg_write_492 = 1'b0 ;
        reg_write_493 = 1'b0 ;
        reg_write_494 = 1'b0 ;
        reg_write_495 = 1'b0 ;
        reg_write_496 = 1'b0 ;
        reg_write_497 = 1'b0 ;
        reg_write_498 = 1'b0 ;
        reg_write_499 = 1'b0 ;
        reg_write_500 = 1'b0 ;
        reg_write_501 = 1'b0 ;
        reg_write_502 = 1'b0 ;
        reg_write_503 = 1'b0 ;
        reg_write_504 = 1'b0 ;
        reg_write_505 = 1'b0 ;
        reg_write_506 = 1'b0 ;
        reg_write_507 = 1'b0 ;
        reg_write_508 = 1'b0 ;
        reg_write_509 = 1'b0 ;
        reg_write_510 = 1'b0 ;
        reg_write_511 = 1'b0 ;
        reg_write_512 = 1'b0 ;
        reg_write_513 = 1'b0 ;
        reg_write_514 = 1'b0 ;
        reg_write_515 = 1'b0 ;
        reg_write_516 = 1'b0 ;
        reg_write_517 = 1'b0 ;
        reg_write_518 = 1'b0 ;
        reg_write_519 = 1'b0 ;
        reg_write_520 = 1'b0 ;
        reg_write_521 = 1'b0 ;
        reg_write_522 = 1'b0 ;
        reg_write_523 = 1'b0 ;
        reg_write_524 = 1'b0 ;
        reg_write_525 = 1'b0 ;
        reg_write_526 = 1'b0 ;
        reg_write_527 = 1'b0 ;
        reg_write_528 = 1'b0 ;
        reg_write_529 = 1'b0 ;
        reg_write_530 = 1'b0 ;
        reg_write_531 = 1'b0 ;
        reg_write_532 = 1'b0 ;
        reg_write_533 = 1'b0 ;
        reg_write_534 = 1'b0 ;
        reg_write_535 = 1'b0 ;
        reg_write_536 = 1'b0 ;
        reg_write_537 = 1'b0 ;
        reg_write_538 = 1'b0 ;
        reg_write_539 = 1'b0 ;
        reg_write_540 = 1'b0 ;
        reg_write_541 = 1'b0 ;
        reg_write_542 = 1'b0 ;
        reg_write_543 = 1'b0 ;
        reg_write_544 = 1'b0 ;
        reg_write_545 = 1'b0 ;
        reg_write_546 = 1'b0 ;
        reg_write_547 = 1'b0 ;
        reg_write_548 = 1'b0 ;
        reg_write_549 = 1'b0 ;
        reg_write_550 = 1'b0 ;
        reg_write_551 = 1'b0 ;
        reg_write_552 = 1'b0 ;
        reg_write_553 = 1'b0 ;
        reg_write_554 = 1'b0 ;
        reg_write_555 = 1'b0 ;
        reg_write_556 = 1'b0 ;
        reg_write_557 = 1'b0 ;
        reg_write_558 = 1'b0 ;
        reg_write_559 = 1'b0 ;
        reg_write_560 = 1'b0 ;
        reg_write_561 = 1'b0 ;
        reg_write_562 = 1'b0 ;
        reg_write_563 = 1'b0 ;
        reg_write_564 = 1'b0 ;
        reg_write_565 = 1'b0 ;
        reg_write_566 = 1'b0 ;
        reg_write_567 = 1'b0 ;
        reg_write_568 = 1'b0 ;
        reg_write_569 = 1'b0 ;
        reg_write_570 = 1'b0 ;
        reg_write_571 = 1'b0 ;
        reg_write_572 = 1'b0 ;
        reg_write_573 = 1'b0 ;
        reg_write_574 = 1'b0 ;
        reg_write_575 = 1'b0 ;
        reg_write_576 = 1'b0 ;
        reg_write_577 = 1'b0 ;
        reg_write_578 = 1'b0 ;
        reg_write_579 = 1'b0 ;
        reg_write_580 = 1'b0 ;
        reg_write_581 = 1'b0 ;
        reg_write_582 = 1'b0 ;
        reg_write_583 = 1'b0 ;
        reg_write_584 = 1'b0 ;
        reg_write_585 = 1'b0 ;
        reg_write_586 = 1'b0 ;
        reg_write_587 = 1'b0 ;
        reg_write_588 = 1'b0 ;
        reg_write_589 = 1'b0 ;
        reg_write_590 = 1'b0 ;
        reg_write_591 = 1'b0 ;
        reg_write_592 = 1'b0 ;
        reg_write_593 = 1'b0 ;
        reg_write_594 = 1'b0 ;
        reg_write_595 = 1'b0 ;
        reg_write_596 = 1'b0 ;
        reg_write_597 = 1'b0 ;
        reg_write_598 = 1'b0 ;
        reg_write_599 = 1'b0 ;
        reg_write_600 = 1'b0 ;
        reg_write_601 = 1'b0 ;
        reg_write_602 = 1'b0 ;
        reg_write_603 = 1'b0 ;
        reg_write_604 = 1'b0 ;
        reg_write_605 = 1'b0 ;
        reg_write_606 = 1'b0 ;
        reg_write_607 = 1'b0 ;
        reg_write_608 = 1'b0 ;
        reg_write_609 = 1'b0 ;
        reg_write_610 = 1'b0 ;
        reg_write_611 = 1'b0 ;
        reg_write_612 = 1'b0 ;
        reg_write_613 = 1'b0 ;
        reg_write_614 = 1'b0 ;
        reg_write_615 = 1'b0 ;
        reg_write_616 = 1'b0 ;
        reg_write_617 = 1'b0 ;
        reg_write_618 = 1'b0 ;
        reg_write_619 = 1'b0 ;
        reg_write_620 = 1'b0 ;
        reg_write_621 = 1'b0 ;
        reg_write_622 = 1'b0 ;
        reg_write_623 = 1'b0 ;
        reg_write_624 = 1'b0 ;
        reg_write_625 = 1'b0 ;
        reg_write_626 = 1'b0 ;
        reg_write_627 = 1'b0 ;
        reg_write_628 = 1'b0 ;
        reg_write_629 = 1'b0 ;
        reg_write_630 = 1'b0 ;
        reg_write_631 = 1'b0 ;
        reg_write_632 = 1'b0 ;
        reg_write_633 = 1'b0 ;
        reg_write_634 = 1'b0 ;
        reg_write_635 = 1'b0 ;
        reg_write_636 = 1'b0 ;
        reg_write_637 = 1'b0 ;
        reg_write_638 = 1'b0 ;
        reg_write_639 = 1'b0 ;
        reg_write_640 = 1'b0 ;
        reg_write_641 = 1'b0 ;
        reg_write_642 = 1'b0 ;
        reg_write_643 = 1'b0 ;
        reg_write_644 = 1'b0 ;
        reg_write_645 = 1'b0 ;
        reg_write_646 = 1'b0 ;
        reg_write_647 = 1'b0 ;
        reg_write_648 = 1'b0 ;
        reg_write_649 = 1'b0 ;
        reg_write_650 = 1'b0 ;
        reg_write_651 = 1'b0 ;
        reg_write_652 = 1'b0 ;
        reg_write_653 = 1'b0 ;
        reg_write_654 = 1'b0 ;
        reg_write_655 = 1'b0 ;
        reg_write_656 = 1'b0 ;
        reg_write_657 = 1'b0 ;
        reg_write_658 = 1'b0 ;
        reg_write_659 = 1'b0 ;
        reg_write_660 = 1'b0 ;
        reg_write_661 = 1'b0 ;
        reg_write_662 = 1'b0 ;
        reg_write_663 = 1'b0 ;
        reg_write_664 = 1'b0 ;
        reg_write_665 = 1'b0 ;
        reg_write_666 = 1'b0 ;
        reg_write_667 = 1'b0 ;
        reg_write_668 = 1'b0 ;
        reg_write_669 = 1'b0 ;
        reg_write_670 = 1'b0 ;
        reg_write_671 = 1'b0 ;
        reg_write_672 = 1'b0 ;
        reg_write_673 = 1'b0 ;
        reg_write_674 = 1'b0 ;
        reg_write_675 = 1'b0 ;
        reg_write_676 = 1'b0 ;
        reg_write_677 = 1'b0 ;
        reg_write_678 = 1'b0 ;
        reg_write_679 = 1'b0 ;
        reg_write_680 = 1'b0 ;
        reg_write_681 = 1'b0 ;
        reg_write_682 = 1'b0 ;
        reg_write_683 = 1'b0 ;
        reg_write_684 = 1'b0 ;
        reg_write_685 = 1'b0 ;
        reg_write_686 = 1'b0 ;
        reg_write_687 = 1'b0 ;
        reg_write_688 = 1'b0 ;
        reg_write_689 = 1'b0 ;
        reg_write_690 = 1'b0 ;
        reg_write_691 = 1'b0 ;
        reg_write_692 = 1'b0 ;
        reg_write_693 = 1'b0 ;
        reg_write_694 = 1'b0 ;
        reg_write_695 = 1'b0 ;
        reg_write_696 = 1'b0 ;
        reg_write_697 = 1'b0 ;
        reg_write_698 = 1'b0 ;
        reg_write_699 = 1'b0 ;
        reg_write_700 = 1'b0 ;
        reg_write_701 = 1'b0 ;
        reg_write_702 = 1'b0 ;
        reg_write_703 = 1'b0 ;
        reg_write_704 = 1'b0 ;
        reg_write_705 = 1'b0 ;
        reg_write_706 = 1'b0 ;
        reg_write_707 = 1'b0 ;
        reg_write_708 = 1'b0 ;
        reg_write_709 = 1'b0 ;
        reg_write_710 = 1'b0 ;
        reg_write_711 = 1'b0 ;
        reg_write_712 = 1'b0 ;
        reg_write_713 = 1'b0 ;
        reg_write_714 = 1'b0 ;
        reg_write_715 = 1'b0 ;
        reg_write_716 = 1'b0 ;
        reg_write_717 = 1'b0 ;
        reg_write_718 = 1'b0 ;
        reg_write_719 = 1'b0 ;
        reg_write_720 = 1'b0 ;
        reg_write_721 = 1'b0 ;
        reg_write_722 = 1'b0 ;
        reg_write_723 = 1'b0 ;
        reg_write_724 = 1'b0 ;
        reg_write_725 = 1'b0 ;
        reg_write_726 = 1'b0 ;
        reg_write_727 = 1'b0 ;
        reg_write_728 = 1'b0 ;
        reg_write_729 = 1'b0 ;
        reg_write_730 = 1'b0 ;
        reg_write_731 = 1'b0 ;
        reg_write_732 = 1'b0 ;
        reg_write_733 = 1'b0 ;
        reg_write_734 = 1'b0 ;
        reg_write_735 = 1'b0 ;
        reg_write_736 = 1'b0 ;
        reg_write_737 = 1'b0 ;
        reg_write_738 = 1'b0 ;
        reg_write_739 = 1'b0 ;
        reg_write_740 = 1'b0 ;
        reg_write_741 = 1'b0 ;
        reg_write_742 = 1'b0 ;
        reg_write_743 = 1'b0 ;
        reg_write_744 = 1'b0 ;
        reg_write_745 = 1'b0 ;
        reg_write_746 = 1'b0 ;
        reg_write_747 = 1'b0 ;
        reg_write_748 = 1'b0 ;
        reg_write_749 = 1'b0 ;
        reg_write_750 = 1'b0 ;
        reg_write_751 = 1'b0 ;
        reg_write_752 = 1'b0 ;
        reg_write_753 = 1'b0 ;
        reg_write_754 = 1'b0 ;
        reg_write_755 = 1'b0 ;
        reg_write_756 = 1'b0 ;
        reg_write_757 = 1'b0 ;
        reg_write_758 = 1'b0 ;
        reg_write_759 = 1'b0 ;
        reg_write_760 = 1'b0 ;
        reg_write_761 = 1'b0 ;
        reg_write_762 = 1'b0 ;
        reg_write_763 = 1'b0 ;
        reg_write_764 = 1'b0 ;
        reg_write_765 = 1'b0 ;
        reg_write_766 = 1'b0 ;
        reg_write_767 = 1'b0 ;
        reg_write_768 = 1'b0 ;
        reg_write_769 = 1'b0 ;
        reg_write_770 = 1'b0 ;
        reg_write_771 = 1'b0 ;
        reg_write_772 = 1'b0 ;
        reg_write_773 = 1'b0 ;
        reg_write_774 = 1'b0 ;
        reg_write_775 = 1'b0 ;
        reg_write_776 = 1'b0 ;
        reg_write_777 = 1'b0 ;
        reg_write_778 = 1'b0 ;
        reg_write_779 = 1'b0 ;
        reg_write_780 = 1'b0 ;
        reg_write_781 = 1'b0 ;
        reg_write_782 = 1'b0 ;
        reg_write_783 = 1'b0 ;
        reg_write_784 = 1'b0 ;
        reg_write_785 = 1'b0 ;
        reg_write_786 = 1'b0 ;
        reg_write_787 = 1'b0 ;
        reg_write_788 = 1'b0 ;
        reg_write_789 = 1'b0 ;
        reg_write_790 = 1'b0 ;
        reg_write_791 = 1'b0 ;
        reg_write_792 = 1'b0 ;
        reg_write_793 = 1'b0 ;
        reg_write_794 = 1'b0 ;
        reg_write_795 = 1'b0 ;
        reg_write_796 = 1'b0 ;
        reg_write_797 = 1'b0 ;
        reg_write_798 = 1'b0 ;
        reg_write_799 = 1'b0 ;
        reg_write_800 = 1'b0 ;
        reg_write_801 = 1'b0 ;
        reg_write_802 = 1'b0 ;
        reg_write_803 = 1'b0 ;
        reg_write_804 = 1'b0 ;
        reg_write_805 = 1'b0 ;
        reg_write_806 = 1'b0 ;
        reg_write_807 = 1'b0 ;
        reg_write_808 = 1'b0 ;
        reg_write_809 = 1'b0 ;
        reg_write_810 = 1'b0 ;
        reg_write_811 = 1'b0 ;
        reg_write_812 = 1'b0 ;
        reg_write_813 = 1'b0 ;
        reg_write_814 = 1'b0 ;
        reg_write_815 = 1'b0 ;
        reg_write_816 = 1'b0 ;
        reg_write_817 = 1'b0 ;
        reg_write_818 = 1'b0 ;
        reg_write_819 = 1'b0 ;
        reg_write_820 = 1'b0 ;
        reg_write_821 = 1'b0 ;
        reg_write_822 = 1'b0 ;
        reg_write_823 = 1'b0 ;
        reg_write_824 = 1'b0 ;
        reg_write_825 = 1'b0 ;
        reg_write_826 = 1'b0 ;
        reg_write_827 = 1'b0 ;
        reg_write_828 = 1'b0 ;
        reg_write_829 = 1'b0 ;
        reg_write_830 = 1'b0 ;
        reg_write_831 = 1'b0 ;
        reg_write_832 = 1'b0 ;
        reg_write_833 = 1'b0 ;
        reg_write_834 = 1'b0 ;
        reg_write_835 = 1'b0 ;
        reg_write_836 = 1'b0 ;
        reg_write_837 = 1'b0 ;
        reg_write_838 = 1'b0 ;
        reg_write_839 = 1'b0 ;
        reg_write_840 = 1'b0 ;
        reg_write_841 = 1'b0 ;
        reg_write_842 = 1'b0 ;
        reg_write_843 = 1'b0 ;
        reg_write_844 = 1'b0 ;
        reg_write_845 = 1'b0 ;
        reg_write_846 = 1'b0 ;
        reg_write_847 = 1'b0 ;
        reg_write_848 = 1'b0 ;
        reg_write_849 = 1'b0 ;
        reg_write_850 = 1'b0 ;
        reg_write_851 = 1'b0 ;
        reg_write_852 = 1'b0 ;
        reg_write_853 = 1'b0 ;
        reg_write_854 = 1'b0 ;
        reg_write_855 = 1'b0 ;
        reg_write_856 = 1'b0 ;
        reg_write_857 = 1'b0 ;
        reg_write_858 = 1'b0 ;
        reg_write_859 = 1'b0 ;
        reg_write_860 = 1'b0 ;
        reg_write_861 = 1'b0 ;
        reg_write_862 = 1'b0 ;
        reg_write_863 = 1'b0 ;
        reg_write_864 = 1'b0 ;
        reg_write_865 = 1'b0 ;
        reg_write_866 = 1'b0 ;
        reg_write_867 = 1'b0 ;
        reg_write_868 = 1'b0 ;
        reg_write_869 = 1'b0 ;
        reg_write_870 = 1'b0 ;
        reg_write_871 = 1'b0 ;
        reg_write_872 = 1'b0 ;
        reg_write_873 = 1'b0 ;
        reg_write_874 = 1'b0 ;
        reg_write_875 = 1'b0 ;
        reg_write_876 = 1'b0 ;
        reg_write_877 = 1'b0 ;
        reg_write_878 = 1'b0 ;
        reg_write_879 = 1'b0 ;
        reg_write_880 = 1'b0 ;
        reg_write_881 = 1'b0 ;
        reg_write_882 = 1'b0 ;
        reg_write_883 = 1'b0 ;
        reg_write_884 = 1'b0 ;
        reg_write_885 = 1'b0 ;
        reg_write_886 = 1'b0 ;
        reg_write_887 = 1'b0 ;
        reg_write_888 = 1'b0 ;
        reg_write_889 = 1'b0 ;
        reg_write_890 = 1'b0 ;
        reg_write_891 = 1'b0 ;
        reg_write_892 = 1'b0 ;
        reg_write_893 = 1'b0 ;
        reg_write_894 = 1'b0 ;
        reg_write_895 = 1'b0 ;
        reg_write_896 = 1'b0 ;
        reg_write_897 = 1'b0 ;
        reg_write_898 = 1'b0 ;
        reg_write_899 = 1'b0 ;
        reg_write_900 = 1'b0 ;
        reg_write_901 = 1'b0 ;
        reg_write_902 = 1'b0 ;
        reg_write_903 = 1'b0 ;
        reg_write_904 = 1'b0 ;
        reg_write_905 = 1'b0 ;
        reg_write_906 = 1'b0 ;
        reg_write_907 = 1'b0 ;
        reg_write_908 = 1'b0 ;
        reg_write_909 = 1'b0 ;
        reg_write_910 = 1'b0 ;
        reg_write_911 = 1'b0 ;
        reg_write_912 = 1'b0 ;
        reg_write_913 = 1'b0 ;
        reg_write_914 = 1'b0 ;
        reg_write_915 = 1'b0 ;
        reg_write_916 = 1'b0 ;
        reg_write_917 = 1'b0 ;
        reg_write_918 = 1'b0 ;
        reg_write_919 = 1'b0 ;
        reg_write_920 = 1'b0 ;
        reg_write_921 = 1'b0 ;
        reg_write_922 = 1'b0 ;
        reg_write_923 = 1'b0 ;
        reg_write_924 = 1'b0 ;
        reg_write_925 = 1'b0 ;
        reg_write_926 = 1'b0 ;
        reg_write_927 = 1'b0 ;
        reg_write_928 = 1'b0 ;
        reg_write_929 = 1'b0 ;
        reg_write_930 = 1'b0 ;
        reg_write_931 = 1'b0 ;
        reg_write_932 = 1'b0 ;
        reg_write_933 = 1'b0 ;
        reg_write_934 = 1'b0 ;
        reg_write_935 = 1'b0 ;
        reg_write_936 = 1'b0 ;
        reg_write_937 = 1'b0 ;
        reg_write_938 = 1'b0 ;
        reg_write_939 = 1'b0 ;
        reg_write_940 = 1'b0 ;
        reg_write_941 = 1'b0 ;
        reg_write_942 = 1'b0 ;
        reg_write_943 = 1'b0 ;
        reg_write_944 = 1'b0 ;
        reg_write_945 = 1'b0 ;
        reg_write_946 = 1'b0 ;
        reg_write_947 = 1'b0 ;
        reg_write_948 = 1'b0 ;
        reg_write_949 = 1'b0 ;
        reg_write_950 = 1'b0 ;
        reg_write_951 = 1'b0 ;
        reg_write_952 = 1'b0 ;
        reg_write_953 = 1'b0 ;
        reg_write_954 = 1'b0 ;
        reg_write_955 = 1'b0 ;
        reg_write_956 = 1'b0 ;
        reg_write_957 = 1'b0 ;
        reg_write_958 = 1'b0 ;
        reg_write_959 = 1'b0 ;
        reg_write_960 = 1'b0 ;
        reg_write_961 = 1'b0 ;
        reg_write_962 = 1'b0 ;
        reg_write_963 = 1'b0 ;
        reg_write_964 = 1'b0 ;
        reg_write_965 = 1'b0 ;
        reg_write_966 = 1'b0 ;
        reg_write_967 = 1'b0 ;
        reg_write_968 = 1'b0 ;
        reg_write_969 = 1'b0 ;
        reg_write_970 = 1'b0 ;
        reg_write_971 = 1'b0 ;
        reg_write_972 = 1'b0 ;
        reg_write_973 = 1'b0 ;
        reg_write_974 = 1'b0 ;
        reg_write_975 = 1'b0 ;
        reg_write_976 = 1'b0 ;
        reg_write_977 = 1'b0 ;
        reg_write_978 = 1'b0 ;
        reg_write_979 = 1'b0 ;
        reg_write_980 = 1'b0 ;
        reg_write_981 = 1'b0 ;
        reg_write_982 = 1'b0 ;
        reg_write_983 = 1'b0 ;
        reg_write_984 = 1'b0 ;
        reg_write_985 = 1'b0 ;
        reg_write_986 = 1'b0 ;
        reg_write_987 = 1'b0 ;
        reg_write_988 = 1'b0 ;
        reg_write_989 = 1'b0 ;
        reg_write_990 = 1'b0 ;
        reg_write_991 = 1'b0 ;
        reg_write_992 = 1'b0 ;
        reg_write_993 = 1'b0 ;
        reg_write_994 = 1'b0 ;
        reg_write_995 = 1'b0 ;
        reg_write_996 = 1'b0 ;
        reg_write_997 = 1'b0 ;
        reg_write_998 = 1'b0 ;
        reg_write_999 = 1'b0 ;
        reg_write_1000 = 1'b0 ;
		if(current_state == 4'd3) begin
			case(counter_ifm) 
        16'd1 : reg_write_1 = 1'b1 ;
        16'd2 : reg_write_2 = 1'b1 ;
        16'd3 : reg_write_3 = 1'b1 ;
        16'd4 : reg_write_4 = 1'b1 ;
        16'd5 : reg_write_5 = 1'b1 ;
        16'd6 : reg_write_6 = 1'b1 ;
        16'd7 : reg_write_7 = 1'b1 ;
        16'd8 : reg_write_8 = 1'b1 ;
        16'd9 : reg_write_9 = 1'b1 ;
        16'd10 : reg_write_10 = 1'b1 ;
        16'd11 : reg_write_11 = 1'b1 ;
        16'd12 : reg_write_12 = 1'b1 ;
        16'd13 : reg_write_13 = 1'b1 ;
        16'd14 : reg_write_14 = 1'b1 ;
        16'd15 : reg_write_15 = 1'b1 ;
        16'd16 : reg_write_16 = 1'b1 ;
        16'd17 : reg_write_17 = 1'b1 ;
        16'd18 : reg_write_18 = 1'b1 ;
        16'd19 : reg_write_19 = 1'b1 ;
        16'd20 : reg_write_20 = 1'b1 ;
        16'd21 : reg_write_21 = 1'b1 ;
        16'd22 : reg_write_22 = 1'b1 ;
        16'd23 : reg_write_23 = 1'b1 ;
        16'd24 : reg_write_24 = 1'b1 ;
        16'd25 : reg_write_25 = 1'b1 ;
        16'd26 : reg_write_26 = 1'b1 ;
        16'd27 : reg_write_27 = 1'b1 ;
        16'd28 : reg_write_28 = 1'b1 ;
        16'd29 : reg_write_29 = 1'b1 ;
        16'd30 : reg_write_30 = 1'b1 ;
        16'd31 : reg_write_31 = 1'b1 ;
        16'd32 : reg_write_32 = 1'b1 ;
        16'd33 : reg_write_33 = 1'b1 ;
        16'd34 : reg_write_34 = 1'b1 ;
        16'd35 : reg_write_35 = 1'b1 ;
        16'd36 : reg_write_36 = 1'b1 ;
        16'd37 : reg_write_37 = 1'b1 ;
        16'd38 : reg_write_38 = 1'b1 ;
        16'd39 : reg_write_39 = 1'b1 ;
        16'd40 : reg_write_40 = 1'b1 ;
        16'd41 : reg_write_41 = 1'b1 ;
        16'd42 : reg_write_42 = 1'b1 ;
        16'd43 : reg_write_43 = 1'b1 ;
        16'd44 : reg_write_44 = 1'b1 ;
        16'd45 : reg_write_45 = 1'b1 ;
        16'd46 : reg_write_46 = 1'b1 ;
        16'd47 : reg_write_47 = 1'b1 ;
        16'd48 : reg_write_48 = 1'b1 ;
        16'd49 : reg_write_49 = 1'b1 ;
        16'd50 : reg_write_50 = 1'b1 ;
        16'd51 : reg_write_51 = 1'b1 ;
        16'd52 : reg_write_52 = 1'b1 ;
        16'd53 : reg_write_53 = 1'b1 ;
        16'd54 : reg_write_54 = 1'b1 ;
        16'd55 : reg_write_55 = 1'b1 ;
        16'd56 : reg_write_56 = 1'b1 ;
        16'd57 : reg_write_57 = 1'b1 ;
        16'd58 : reg_write_58 = 1'b1 ;
        16'd59 : reg_write_59 = 1'b1 ;
        16'd60 : reg_write_60 = 1'b1 ;
        16'd61 : reg_write_61 = 1'b1 ;
        16'd62 : reg_write_62 = 1'b1 ;
        16'd63 : reg_write_63 = 1'b1 ;
        16'd64 : reg_write_64 = 1'b1 ;
        16'd65 : reg_write_65 = 1'b1 ;
        16'd66 : reg_write_66 = 1'b1 ;
        16'd67 : reg_write_67 = 1'b1 ;
        16'd68 : reg_write_68 = 1'b1 ;
        16'd69 : reg_write_69 = 1'b1 ;
        16'd70 : reg_write_70 = 1'b1 ;
        16'd71 : reg_write_71 = 1'b1 ;
        16'd72 : reg_write_72 = 1'b1 ;
        16'd73 : reg_write_73 = 1'b1 ;
        16'd74 : reg_write_74 = 1'b1 ;
        16'd75 : reg_write_75 = 1'b1 ;
        16'd76 : reg_write_76 = 1'b1 ;
        16'd77 : reg_write_77 = 1'b1 ;
        16'd78 : reg_write_78 = 1'b1 ;
        16'd79 : reg_write_79 = 1'b1 ;
        16'd80 : reg_write_80 = 1'b1 ;
        16'd81 : reg_write_81 = 1'b1 ;
        16'd82 : reg_write_82 = 1'b1 ;
        16'd83 : reg_write_83 = 1'b1 ;
        16'd84 : reg_write_84 = 1'b1 ;
        16'd85 : reg_write_85 = 1'b1 ;
        16'd86 : reg_write_86 = 1'b1 ;
        16'd87 : reg_write_87 = 1'b1 ;
        16'd88 : reg_write_88 = 1'b1 ;
        16'd89 : reg_write_89 = 1'b1 ;
        16'd90 : reg_write_90 = 1'b1 ;
        16'd91 : reg_write_91 = 1'b1 ;
        16'd92 : reg_write_92 = 1'b1 ;
        16'd93 : reg_write_93 = 1'b1 ;
        16'd94 : reg_write_94 = 1'b1 ;
        16'd95 : reg_write_95 = 1'b1 ;
        16'd96 : reg_write_96 = 1'b1 ;
        16'd97 : reg_write_97 = 1'b1 ;
        16'd98 : reg_write_98 = 1'b1 ;
        16'd99 : reg_write_99 = 1'b1 ;
        16'd100 : reg_write_100 = 1'b1 ;
        16'd101 : reg_write_101 = 1'b1 ;
        16'd102 : reg_write_102 = 1'b1 ;
        16'd103 : reg_write_103 = 1'b1 ;
        16'd104 : reg_write_104 = 1'b1 ;
        16'd105 : reg_write_105 = 1'b1 ;
        16'd106 : reg_write_106 = 1'b1 ;
        16'd107 : reg_write_107 = 1'b1 ;
        16'd108 : reg_write_108 = 1'b1 ;
        16'd109 : reg_write_109 = 1'b1 ;
        16'd110 : reg_write_110 = 1'b1 ;
        16'd111 : reg_write_111 = 1'b1 ;
        16'd112 : reg_write_112 = 1'b1 ;
        16'd113 : reg_write_113 = 1'b1 ;
        16'd114 : reg_write_114 = 1'b1 ;
        16'd115 : reg_write_115 = 1'b1 ;
        16'd116 : reg_write_116 = 1'b1 ;
        16'd117 : reg_write_117 = 1'b1 ;
        16'd118 : reg_write_118 = 1'b1 ;
        16'd119 : reg_write_119 = 1'b1 ;
        16'd120 : reg_write_120 = 1'b1 ;
        16'd121 : reg_write_121 = 1'b1 ;
        16'd122 : reg_write_122 = 1'b1 ;
        16'd123 : reg_write_123 = 1'b1 ;
        16'd124 : reg_write_124 = 1'b1 ;
        16'd125 : reg_write_125 = 1'b1 ;
        16'd126 : reg_write_126 = 1'b1 ;
        16'd127 : reg_write_127 = 1'b1 ;
        16'd128 : reg_write_128 = 1'b1 ;
        16'd129 : reg_write_129 = 1'b1 ;
        16'd130 : reg_write_130 = 1'b1 ;
        16'd131 : reg_write_131 = 1'b1 ;
        16'd132 : reg_write_132 = 1'b1 ;
        16'd133 : reg_write_133 = 1'b1 ;
        16'd134 : reg_write_134 = 1'b1 ;
        16'd135 : reg_write_135 = 1'b1 ;
        16'd136 : reg_write_136 = 1'b1 ;
        16'd137 : reg_write_137 = 1'b1 ;
        16'd138 : reg_write_138 = 1'b1 ;
        16'd139 : reg_write_139 = 1'b1 ;
        16'd140 : reg_write_140 = 1'b1 ;
        16'd141 : reg_write_141 = 1'b1 ;
        16'd142 : reg_write_142 = 1'b1 ;
        16'd143 : reg_write_143 = 1'b1 ;
        16'd144 : reg_write_144 = 1'b1 ;
        16'd145 : reg_write_145 = 1'b1 ;
        16'd146 : reg_write_146 = 1'b1 ;
        16'd147 : reg_write_147 = 1'b1 ;
        16'd148 : reg_write_148 = 1'b1 ;
        16'd149 : reg_write_149 = 1'b1 ;
        16'd150 : reg_write_150 = 1'b1 ;
        16'd151 : reg_write_151 = 1'b1 ;
        16'd152 : reg_write_152 = 1'b1 ;
        16'd153 : reg_write_153 = 1'b1 ;
        16'd154 : reg_write_154 = 1'b1 ;
        16'd155 : reg_write_155 = 1'b1 ;
        16'd156 : reg_write_156 = 1'b1 ;
        16'd157 : reg_write_157 = 1'b1 ;
        16'd158 : reg_write_158 = 1'b1 ;
        16'd159 : reg_write_159 = 1'b1 ;
        16'd160 : reg_write_160 = 1'b1 ;
        16'd161 : reg_write_161 = 1'b1 ;
        16'd162 : reg_write_162 = 1'b1 ;
        16'd163 : reg_write_163 = 1'b1 ;
        16'd164 : reg_write_164 = 1'b1 ;
        16'd165 : reg_write_165 = 1'b1 ;
        16'd166 : reg_write_166 = 1'b1 ;
        16'd167 : reg_write_167 = 1'b1 ;
        16'd168 : reg_write_168 = 1'b1 ;
        16'd169 : reg_write_169 = 1'b1 ;
        16'd170 : reg_write_170 = 1'b1 ;
        16'd171 : reg_write_171 = 1'b1 ;
        16'd172 : reg_write_172 = 1'b1 ;
        16'd173 : reg_write_173 = 1'b1 ;
        16'd174 : reg_write_174 = 1'b1 ;
        16'd175 : reg_write_175 = 1'b1 ;
        16'd176 : reg_write_176 = 1'b1 ;
        16'd177 : reg_write_177 = 1'b1 ;
        16'd178 : reg_write_178 = 1'b1 ;
        16'd179 : reg_write_179 = 1'b1 ;
        16'd180 : reg_write_180 = 1'b1 ;
        16'd181 : reg_write_181 = 1'b1 ;
        16'd182 : reg_write_182 = 1'b1 ;
        16'd183 : reg_write_183 = 1'b1 ;
        16'd184 : reg_write_184 = 1'b1 ;
        16'd185 : reg_write_185 = 1'b1 ;
        16'd186 : reg_write_186 = 1'b1 ;
        16'd187 : reg_write_187 = 1'b1 ;
        16'd188 : reg_write_188 = 1'b1 ;
        16'd189 : reg_write_189 = 1'b1 ;
        16'd190 : reg_write_190 = 1'b1 ;
        16'd191 : reg_write_191 = 1'b1 ;
        16'd192 : reg_write_192 = 1'b1 ;
        16'd193 : reg_write_193 = 1'b1 ;
        16'd194 : reg_write_194 = 1'b1 ;
        16'd195 : reg_write_195 = 1'b1 ;
        16'd196 : reg_write_196 = 1'b1 ;
        16'd197 : reg_write_197 = 1'b1 ;
        16'd198 : reg_write_198 = 1'b1 ;
        16'd199 : reg_write_199 = 1'b1 ;
        16'd200 : reg_write_200 = 1'b1 ;
        16'd201 : reg_write_201 = 1'b1 ;
        16'd202 : reg_write_202 = 1'b1 ;
        16'd203 : reg_write_203 = 1'b1 ;
        16'd204 : reg_write_204 = 1'b1 ;
        16'd205 : reg_write_205 = 1'b1 ;
        16'd206 : reg_write_206 = 1'b1 ;
        16'd207 : reg_write_207 = 1'b1 ;
        16'd208 : reg_write_208 = 1'b1 ;
        16'd209 : reg_write_209 = 1'b1 ;
        16'd210 : reg_write_210 = 1'b1 ;
        16'd211 : reg_write_211 = 1'b1 ;
        16'd212 : reg_write_212 = 1'b1 ;
        16'd213 : reg_write_213 = 1'b1 ;
        16'd214 : reg_write_214 = 1'b1 ;
        16'd215 : reg_write_215 = 1'b1 ;
        16'd216 : reg_write_216 = 1'b1 ;
        16'd217 : reg_write_217 = 1'b1 ;
        16'd218 : reg_write_218 = 1'b1 ;
        16'd219 : reg_write_219 = 1'b1 ;
        16'd220 : reg_write_220 = 1'b1 ;
        16'd221 : reg_write_221 = 1'b1 ;
        16'd222 : reg_write_222 = 1'b1 ;
        16'd223 : reg_write_223 = 1'b1 ;
        16'd224 : reg_write_224 = 1'b1 ;
        16'd225 : reg_write_225 = 1'b1 ;
        16'd226 : reg_write_226 = 1'b1 ;
        16'd227 : reg_write_227 = 1'b1 ;
        16'd228 : reg_write_228 = 1'b1 ;
        16'd229 : reg_write_229 = 1'b1 ;
        16'd230 : reg_write_230 = 1'b1 ;
        16'd231 : reg_write_231 = 1'b1 ;
        16'd232 : reg_write_232 = 1'b1 ;
        16'd233 : reg_write_233 = 1'b1 ;
        16'd234 : reg_write_234 = 1'b1 ;
        16'd235 : reg_write_235 = 1'b1 ;
        16'd236 : reg_write_236 = 1'b1 ;
        16'd237 : reg_write_237 = 1'b1 ;
        16'd238 : reg_write_238 = 1'b1 ;
        16'd239 : reg_write_239 = 1'b1 ;
        16'd240 : reg_write_240 = 1'b1 ;
        16'd241 : reg_write_241 = 1'b1 ;
        16'd242 : reg_write_242 = 1'b1 ;
        16'd243 : reg_write_243 = 1'b1 ;
        16'd244 : reg_write_244 = 1'b1 ;
        16'd245 : reg_write_245 = 1'b1 ;
        16'd246 : reg_write_246 = 1'b1 ;
        16'd247 : reg_write_247 = 1'b1 ;
        16'd248 : reg_write_248 = 1'b1 ;
        16'd249 : reg_write_249 = 1'b1 ;
        16'd250 : reg_write_250 = 1'b1 ;
        16'd251 : reg_write_251 = 1'b1 ;
        16'd252 : reg_write_252 = 1'b1 ;
        16'd253 : reg_write_253 = 1'b1 ;
        16'd254 : reg_write_254 = 1'b1 ;
        16'd255 : reg_write_255 = 1'b1 ;
        16'd256 : reg_write_256 = 1'b1 ;
        16'd257 : reg_write_257 = 1'b1 ;
        16'd258 : reg_write_258 = 1'b1 ;
        16'd259 : reg_write_259 = 1'b1 ;
        16'd260 : reg_write_260 = 1'b1 ;
        16'd261 : reg_write_261 = 1'b1 ;
        16'd262 : reg_write_262 = 1'b1 ;
        16'd263 : reg_write_263 = 1'b1 ;
        16'd264 : reg_write_264 = 1'b1 ;
        16'd265 : reg_write_265 = 1'b1 ;
        16'd266 : reg_write_266 = 1'b1 ;
        16'd267 : reg_write_267 = 1'b1 ;
        16'd268 : reg_write_268 = 1'b1 ;
        16'd269 : reg_write_269 = 1'b1 ;
        16'd270 : reg_write_270 = 1'b1 ;
        16'd271 : reg_write_271 = 1'b1 ;
        16'd272 : reg_write_272 = 1'b1 ;
        16'd273 : reg_write_273 = 1'b1 ;
        16'd274 : reg_write_274 = 1'b1 ;
        16'd275 : reg_write_275 = 1'b1 ;
        16'd276 : reg_write_276 = 1'b1 ;
        16'd277 : reg_write_277 = 1'b1 ;
        16'd278 : reg_write_278 = 1'b1 ;
        16'd279 : reg_write_279 = 1'b1 ;
        16'd280 : reg_write_280 = 1'b1 ;
        16'd281 : reg_write_281 = 1'b1 ;
        16'd282 : reg_write_282 = 1'b1 ;
        16'd283 : reg_write_283 = 1'b1 ;
        16'd284 : reg_write_284 = 1'b1 ;
        16'd285 : reg_write_285 = 1'b1 ;
        16'd286 : reg_write_286 = 1'b1 ;
        16'd287 : reg_write_287 = 1'b1 ;
        16'd288 : reg_write_288 = 1'b1 ;
        16'd289 : reg_write_289 = 1'b1 ;
        16'd290 : reg_write_290 = 1'b1 ;
        16'd291 : reg_write_291 = 1'b1 ;
        16'd292 : reg_write_292 = 1'b1 ;
        16'd293 : reg_write_293 = 1'b1 ;
        16'd294 : reg_write_294 = 1'b1 ;
        16'd295 : reg_write_295 = 1'b1 ;
        16'd296 : reg_write_296 = 1'b1 ;
        16'd297 : reg_write_297 = 1'b1 ;
        16'd298 : reg_write_298 = 1'b1 ;
        16'd299 : reg_write_299 = 1'b1 ;
        16'd300 : reg_write_300 = 1'b1 ;
        16'd301 : reg_write_301 = 1'b1 ;
        16'd302 : reg_write_302 = 1'b1 ;
        16'd303 : reg_write_303 = 1'b1 ;
        16'd304 : reg_write_304 = 1'b1 ;
        16'd305 : reg_write_305 = 1'b1 ;
        16'd306 : reg_write_306 = 1'b1 ;
        16'd307 : reg_write_307 = 1'b1 ;
        16'd308 : reg_write_308 = 1'b1 ;
        16'd309 : reg_write_309 = 1'b1 ;
        16'd310 : reg_write_310 = 1'b1 ;
        16'd311 : reg_write_311 = 1'b1 ;
        16'd312 : reg_write_312 = 1'b1 ;
        16'd313 : reg_write_313 = 1'b1 ;
        16'd314 : reg_write_314 = 1'b1 ;
        16'd315 : reg_write_315 = 1'b1 ;
        16'd316 : reg_write_316 = 1'b1 ;
        16'd317 : reg_write_317 = 1'b1 ;
        16'd318 : reg_write_318 = 1'b1 ;
        16'd319 : reg_write_319 = 1'b1 ;
        16'd320 : reg_write_320 = 1'b1 ;
        16'd321 : reg_write_321 = 1'b1 ;
        16'd322 : reg_write_322 = 1'b1 ;
        16'd323 : reg_write_323 = 1'b1 ;
        16'd324 : reg_write_324 = 1'b1 ;
        16'd325 : reg_write_325 = 1'b1 ;
        16'd326 : reg_write_326 = 1'b1 ;
        16'd327 : reg_write_327 = 1'b1 ;
        16'd328 : reg_write_328 = 1'b1 ;
        16'd329 : reg_write_329 = 1'b1 ;
        16'd330 : reg_write_330 = 1'b1 ;
        16'd331 : reg_write_331 = 1'b1 ;
        16'd332 : reg_write_332 = 1'b1 ;
        16'd333 : reg_write_333 = 1'b1 ;
        16'd334 : reg_write_334 = 1'b1 ;
        16'd335 : reg_write_335 = 1'b1 ;
        16'd336 : reg_write_336 = 1'b1 ;
        16'd337 : reg_write_337 = 1'b1 ;
        16'd338 : reg_write_338 = 1'b1 ;
        16'd339 : reg_write_339 = 1'b1 ;
        16'd340 : reg_write_340 = 1'b1 ;
        16'd341 : reg_write_341 = 1'b1 ;
        16'd342 : reg_write_342 = 1'b1 ;
        16'd343 : reg_write_343 = 1'b1 ;
        16'd344 : reg_write_344 = 1'b1 ;
        16'd345 : reg_write_345 = 1'b1 ;
        16'd346 : reg_write_346 = 1'b1 ;
        16'd347 : reg_write_347 = 1'b1 ;
        16'd348 : reg_write_348 = 1'b1 ;
        16'd349 : reg_write_349 = 1'b1 ;
        16'd350 : reg_write_350 = 1'b1 ;
        16'd351 : reg_write_351 = 1'b1 ;
        16'd352 : reg_write_352 = 1'b1 ;
        16'd353 : reg_write_353 = 1'b1 ;
        16'd354 : reg_write_354 = 1'b1 ;
        16'd355 : reg_write_355 = 1'b1 ;
        16'd356 : reg_write_356 = 1'b1 ;
        16'd357 : reg_write_357 = 1'b1 ;
        16'd358 : reg_write_358 = 1'b1 ;
        16'd359 : reg_write_359 = 1'b1 ;
        16'd360 : reg_write_360 = 1'b1 ;
        16'd361 : reg_write_361 = 1'b1 ;
        16'd362 : reg_write_362 = 1'b1 ;
        16'd363 : reg_write_363 = 1'b1 ;
        16'd364 : reg_write_364 = 1'b1 ;
        16'd365 : reg_write_365 = 1'b1 ;
        16'd366 : reg_write_366 = 1'b1 ;
        16'd367 : reg_write_367 = 1'b1 ;
        16'd368 : reg_write_368 = 1'b1 ;
        16'd369 : reg_write_369 = 1'b1 ;
        16'd370 : reg_write_370 = 1'b1 ;
        16'd371 : reg_write_371 = 1'b1 ;
        16'd372 : reg_write_372 = 1'b1 ;
        16'd373 : reg_write_373 = 1'b1 ;
        16'd374 : reg_write_374 = 1'b1 ;
        16'd375 : reg_write_375 = 1'b1 ;
        16'd376 : reg_write_376 = 1'b1 ;
        16'd377 : reg_write_377 = 1'b1 ;
        16'd378 : reg_write_378 = 1'b1 ;
        16'd379 : reg_write_379 = 1'b1 ;
        16'd380 : reg_write_380 = 1'b1 ;
        16'd381 : reg_write_381 = 1'b1 ;
        16'd382 : reg_write_382 = 1'b1 ;
        16'd383 : reg_write_383 = 1'b1 ;
        16'd384 : reg_write_384 = 1'b1 ;
        16'd385 : reg_write_385 = 1'b1 ;
        16'd386 : reg_write_386 = 1'b1 ;
        16'd387 : reg_write_387 = 1'b1 ;
        16'd388 : reg_write_388 = 1'b1 ;
        16'd389 : reg_write_389 = 1'b1 ;
        16'd390 : reg_write_390 = 1'b1 ;
        16'd391 : reg_write_391 = 1'b1 ;
        16'd392 : reg_write_392 = 1'b1 ;
        16'd393 : reg_write_393 = 1'b1 ;
        16'd394 : reg_write_394 = 1'b1 ;
        16'd395 : reg_write_395 = 1'b1 ;
        16'd396 : reg_write_396 = 1'b1 ;
        16'd397 : reg_write_397 = 1'b1 ;
        16'd398 : reg_write_398 = 1'b1 ;
        16'd399 : reg_write_399 = 1'b1 ;
        16'd400 : reg_write_400 = 1'b1 ;
        16'd401 : reg_write_401 = 1'b1 ;
        16'd402 : reg_write_402 = 1'b1 ;
        16'd403 : reg_write_403 = 1'b1 ;
        16'd404 : reg_write_404 = 1'b1 ;
        16'd405 : reg_write_405 = 1'b1 ;
        16'd406 : reg_write_406 = 1'b1 ;
        16'd407 : reg_write_407 = 1'b1 ;
        16'd408 : reg_write_408 = 1'b1 ;
        16'd409 : reg_write_409 = 1'b1 ;
        16'd410 : reg_write_410 = 1'b1 ;
        16'd411 : reg_write_411 = 1'b1 ;
        16'd412 : reg_write_412 = 1'b1 ;
        16'd413 : reg_write_413 = 1'b1 ;
        16'd414 : reg_write_414 = 1'b1 ;
        16'd415 : reg_write_415 = 1'b1 ;
        16'd416 : reg_write_416 = 1'b1 ;
        16'd417 : reg_write_417 = 1'b1 ;
        16'd418 : reg_write_418 = 1'b1 ;
        16'd419 : reg_write_419 = 1'b1 ;
        16'd420 : reg_write_420 = 1'b1 ;
        16'd421 : reg_write_421 = 1'b1 ;
        16'd422 : reg_write_422 = 1'b1 ;
        16'd423 : reg_write_423 = 1'b1 ;
        16'd424 : reg_write_424 = 1'b1 ;
        16'd425 : reg_write_425 = 1'b1 ;
        16'd426 : reg_write_426 = 1'b1 ;
        16'd427 : reg_write_427 = 1'b1 ;
        16'd428 : reg_write_428 = 1'b1 ;
        16'd429 : reg_write_429 = 1'b1 ;
        16'd430 : reg_write_430 = 1'b1 ;
        16'd431 : reg_write_431 = 1'b1 ;
        16'd432 : reg_write_432 = 1'b1 ;
        16'd433 : reg_write_433 = 1'b1 ;
        16'd434 : reg_write_434 = 1'b1 ;
        16'd435 : reg_write_435 = 1'b1 ;
        16'd436 : reg_write_436 = 1'b1 ;
        16'd437 : reg_write_437 = 1'b1 ;
        16'd438 : reg_write_438 = 1'b1 ;
        16'd439 : reg_write_439 = 1'b1 ;
        16'd440 : reg_write_440 = 1'b1 ;
        16'd441 : reg_write_441 = 1'b1 ;
        16'd442 : reg_write_442 = 1'b1 ;
        16'd443 : reg_write_443 = 1'b1 ;
        16'd444 : reg_write_444 = 1'b1 ;
        16'd445 : reg_write_445 = 1'b1 ;
        16'd446 : reg_write_446 = 1'b1 ;
        16'd447 : reg_write_447 = 1'b1 ;
        16'd448 : reg_write_448 = 1'b1 ;
        16'd449 : reg_write_449 = 1'b1 ;
        16'd450 : reg_write_450 = 1'b1 ;
        16'd451 : reg_write_451 = 1'b1 ;
        16'd452 : reg_write_452 = 1'b1 ;
        16'd453 : reg_write_453 = 1'b1 ;
        16'd454 : reg_write_454 = 1'b1 ;
        16'd455 : reg_write_455 = 1'b1 ;
        16'd456 : reg_write_456 = 1'b1 ;
        16'd457 : reg_write_457 = 1'b1 ;
        16'd458 : reg_write_458 = 1'b1 ;
        16'd459 : reg_write_459 = 1'b1 ;
        16'd460 : reg_write_460 = 1'b1 ;
        16'd461 : reg_write_461 = 1'b1 ;
        16'd462 : reg_write_462 = 1'b1 ;
        16'd463 : reg_write_463 = 1'b1 ;
        16'd464 : reg_write_464 = 1'b1 ;
        16'd465 : reg_write_465 = 1'b1 ;
        16'd466 : reg_write_466 = 1'b1 ;
        16'd467 : reg_write_467 = 1'b1 ;
        16'd468 : reg_write_468 = 1'b1 ;
        16'd469 : reg_write_469 = 1'b1 ;
        16'd470 : reg_write_470 = 1'b1 ;
        16'd471 : reg_write_471 = 1'b1 ;
        16'd472 : reg_write_472 = 1'b1 ;
        16'd473 : reg_write_473 = 1'b1 ;
        16'd474 : reg_write_474 = 1'b1 ;
        16'd475 : reg_write_475 = 1'b1 ;
        16'd476 : reg_write_476 = 1'b1 ;
        16'd477 : reg_write_477 = 1'b1 ;
        16'd478 : reg_write_478 = 1'b1 ;
        16'd479 : reg_write_479 = 1'b1 ;
        16'd480 : reg_write_480 = 1'b1 ;
        16'd481 : reg_write_481 = 1'b1 ;
        16'd482 : reg_write_482 = 1'b1 ;
        16'd483 : reg_write_483 = 1'b1 ;
        16'd484 : reg_write_484 = 1'b1 ;
        16'd485 : reg_write_485 = 1'b1 ;
        16'd486 : reg_write_486 = 1'b1 ;
        16'd487 : reg_write_487 = 1'b1 ;
        16'd488 : reg_write_488 = 1'b1 ;
        16'd489 : reg_write_489 = 1'b1 ;
        16'd490 : reg_write_490 = 1'b1 ;
        16'd491 : reg_write_491 = 1'b1 ;
        16'd492 : reg_write_492 = 1'b1 ;
        16'd493 : reg_write_493 = 1'b1 ;
        16'd494 : reg_write_494 = 1'b1 ;
        16'd495 : reg_write_495 = 1'b1 ;
        16'd496 : reg_write_496 = 1'b1 ;
        16'd497 : reg_write_497 = 1'b1 ;
        16'd498 : reg_write_498 = 1'b1 ;
        16'd499 : reg_write_499 = 1'b1 ;
        16'd500 : reg_write_500 = 1'b1 ;
        16'd501 : reg_write_501 = 1'b1 ;
        16'd502 : reg_write_502 = 1'b1 ;
        16'd503 : reg_write_503 = 1'b1 ;
        16'd504 : reg_write_504 = 1'b1 ;
        16'd505 : reg_write_505 = 1'b1 ;
        16'd506 : reg_write_506 = 1'b1 ;
        16'd507 : reg_write_507 = 1'b1 ;
        16'd508 : reg_write_508 = 1'b1 ;
        16'd509 : reg_write_509 = 1'b1 ;
        16'd510 : reg_write_510 = 1'b1 ;
        16'd511 : reg_write_511 = 1'b1 ;
        16'd512 : reg_write_512 = 1'b1 ;
        16'd513 : reg_write_513 = 1'b1 ;
        16'd514 : reg_write_514 = 1'b1 ;
        16'd515 : reg_write_515 = 1'b1 ;
        16'd516 : reg_write_516 = 1'b1 ;
        16'd517 : reg_write_517 = 1'b1 ;
        16'd518 : reg_write_518 = 1'b1 ;
        16'd519 : reg_write_519 = 1'b1 ;
        16'd520 : reg_write_520 = 1'b1 ;
        16'd521 : reg_write_521 = 1'b1 ;
        16'd522 : reg_write_522 = 1'b1 ;
        16'd523 : reg_write_523 = 1'b1 ;
        16'd524 : reg_write_524 = 1'b1 ;
        16'd525 : reg_write_525 = 1'b1 ;
        16'd526 : reg_write_526 = 1'b1 ;
        16'd527 : reg_write_527 = 1'b1 ;
        16'd528 : reg_write_528 = 1'b1 ;
        16'd529 : reg_write_529 = 1'b1 ;
        16'd530 : reg_write_530 = 1'b1 ;
        16'd531 : reg_write_531 = 1'b1 ;
        16'd532 : reg_write_532 = 1'b1 ;
        16'd533 : reg_write_533 = 1'b1 ;
        16'd534 : reg_write_534 = 1'b1 ;
        16'd535 : reg_write_535 = 1'b1 ;
        16'd536 : reg_write_536 = 1'b1 ;
        16'd537 : reg_write_537 = 1'b1 ;
        16'd538 : reg_write_538 = 1'b1 ;
        16'd539 : reg_write_539 = 1'b1 ;
        16'd540 : reg_write_540 = 1'b1 ;
        16'd541 : reg_write_541 = 1'b1 ;
        16'd542 : reg_write_542 = 1'b1 ;
        16'd543 : reg_write_543 = 1'b1 ;
        16'd544 : reg_write_544 = 1'b1 ;
        16'd545 : reg_write_545 = 1'b1 ;
        16'd546 : reg_write_546 = 1'b1 ;
        16'd547 : reg_write_547 = 1'b1 ;
        16'd548 : reg_write_548 = 1'b1 ;
        16'd549 : reg_write_549 = 1'b1 ;
        16'd550 : reg_write_550 = 1'b1 ;
        16'd551 : reg_write_551 = 1'b1 ;
        16'd552 : reg_write_552 = 1'b1 ;
        16'd553 : reg_write_553 = 1'b1 ;
        16'd554 : reg_write_554 = 1'b1 ;
        16'd555 : reg_write_555 = 1'b1 ;
        16'd556 : reg_write_556 = 1'b1 ;
        16'd557 : reg_write_557 = 1'b1 ;
        16'd558 : reg_write_558 = 1'b1 ;
        16'd559 : reg_write_559 = 1'b1 ;
        16'd560 : reg_write_560 = 1'b1 ;
        16'd561 : reg_write_561 = 1'b1 ;
        16'd562 : reg_write_562 = 1'b1 ;
        16'd563 : reg_write_563 = 1'b1 ;
        16'd564 : reg_write_564 = 1'b1 ;
        16'd565 : reg_write_565 = 1'b1 ;
        16'd566 : reg_write_566 = 1'b1 ;
        16'd567 : reg_write_567 = 1'b1 ;
        16'd568 : reg_write_568 = 1'b1 ;
        16'd569 : reg_write_569 = 1'b1 ;
        16'd570 : reg_write_570 = 1'b1 ;
        16'd571 : reg_write_571 = 1'b1 ;
        16'd572 : reg_write_572 = 1'b1 ;
        16'd573 : reg_write_573 = 1'b1 ;
        16'd574 : reg_write_574 = 1'b1 ;
        16'd575 : reg_write_575 = 1'b1 ;
        16'd576 : reg_write_576 = 1'b1 ;
        16'd577 : reg_write_577 = 1'b1 ;
        16'd578 : reg_write_578 = 1'b1 ;
        16'd579 : reg_write_579 = 1'b1 ;
        16'd580 : reg_write_580 = 1'b1 ;
        16'd581 : reg_write_581 = 1'b1 ;
        16'd582 : reg_write_582 = 1'b1 ;
        16'd583 : reg_write_583 = 1'b1 ;
        16'd584 : reg_write_584 = 1'b1 ;
        16'd585 : reg_write_585 = 1'b1 ;
        16'd586 : reg_write_586 = 1'b1 ;
        16'd587 : reg_write_587 = 1'b1 ;
        16'd588 : reg_write_588 = 1'b1 ;
        16'd589 : reg_write_589 = 1'b1 ;
        16'd590 : reg_write_590 = 1'b1 ;
        16'd591 : reg_write_591 = 1'b1 ;
        16'd592 : reg_write_592 = 1'b1 ;
        16'd593 : reg_write_593 = 1'b1 ;
        16'd594 : reg_write_594 = 1'b1 ;
        16'd595 : reg_write_595 = 1'b1 ;
        16'd596 : reg_write_596 = 1'b1 ;
        16'd597 : reg_write_597 = 1'b1 ;
        16'd598 : reg_write_598 = 1'b1 ;
        16'd599 : reg_write_599 = 1'b1 ;
        16'd600 : reg_write_600 = 1'b1 ;
        16'd601 : reg_write_601 = 1'b1 ;
        16'd602 : reg_write_602 = 1'b1 ;
        16'd603 : reg_write_603 = 1'b1 ;
        16'd604 : reg_write_604 = 1'b1 ;
        16'd605 : reg_write_605 = 1'b1 ;
        16'd606 : reg_write_606 = 1'b1 ;
        16'd607 : reg_write_607 = 1'b1 ;
        16'd608 : reg_write_608 = 1'b1 ;
        16'd609 : reg_write_609 = 1'b1 ;
        16'd610 : reg_write_610 = 1'b1 ;
        16'd611 : reg_write_611 = 1'b1 ;
        16'd612 : reg_write_612 = 1'b1 ;
        16'd613 : reg_write_613 = 1'b1 ;
        16'd614 : reg_write_614 = 1'b1 ;
        16'd615 : reg_write_615 = 1'b1 ;
        16'd616 : reg_write_616 = 1'b1 ;
        16'd617 : reg_write_617 = 1'b1 ;
        16'd618 : reg_write_618 = 1'b1 ;
        16'd619 : reg_write_619 = 1'b1 ;
        16'd620 : reg_write_620 = 1'b1 ;
        16'd621 : reg_write_621 = 1'b1 ;
        16'd622 : reg_write_622 = 1'b1 ;
        16'd623 : reg_write_623 = 1'b1 ;
        16'd624 : reg_write_624 = 1'b1 ;
        16'd625 : reg_write_625 = 1'b1 ;
        16'd626 : reg_write_626 = 1'b1 ;
        16'd627 : reg_write_627 = 1'b1 ;
        16'd628 : reg_write_628 = 1'b1 ;
        16'd629 : reg_write_629 = 1'b1 ;
        16'd630 : reg_write_630 = 1'b1 ;
        16'd631 : reg_write_631 = 1'b1 ;
        16'd632 : reg_write_632 = 1'b1 ;
        16'd633 : reg_write_633 = 1'b1 ;
        16'd634 : reg_write_634 = 1'b1 ;
        16'd635 : reg_write_635 = 1'b1 ;
        16'd636 : reg_write_636 = 1'b1 ;
        16'd637 : reg_write_637 = 1'b1 ;
        16'd638 : reg_write_638 = 1'b1 ;
        16'd639 : reg_write_639 = 1'b1 ;
        16'd640 : reg_write_640 = 1'b1 ;
        16'd641 : reg_write_641 = 1'b1 ;
        16'd642 : reg_write_642 = 1'b1 ;
        16'd643 : reg_write_643 = 1'b1 ;
        16'd644 : reg_write_644 = 1'b1 ;
        16'd645 : reg_write_645 = 1'b1 ;
        16'd646 : reg_write_646 = 1'b1 ;
        16'd647 : reg_write_647 = 1'b1 ;
        16'd648 : reg_write_648 = 1'b1 ;
        16'd649 : reg_write_649 = 1'b1 ;
        16'd650 : reg_write_650 = 1'b1 ;
        16'd651 : reg_write_651 = 1'b1 ;
        16'd652 : reg_write_652 = 1'b1 ;
        16'd653 : reg_write_653 = 1'b1 ;
        16'd654 : reg_write_654 = 1'b1 ;
        16'd655 : reg_write_655 = 1'b1 ;
        16'd656 : reg_write_656 = 1'b1 ;
        16'd657 : reg_write_657 = 1'b1 ;
        16'd658 : reg_write_658 = 1'b1 ;
        16'd659 : reg_write_659 = 1'b1 ;
        16'd660 : reg_write_660 = 1'b1 ;
        16'd661 : reg_write_661 = 1'b1 ;
        16'd662 : reg_write_662 = 1'b1 ;
        16'd663 : reg_write_663 = 1'b1 ;
        16'd664 : reg_write_664 = 1'b1 ;
        16'd665 : reg_write_665 = 1'b1 ;
        16'd666 : reg_write_666 = 1'b1 ;
        16'd667 : reg_write_667 = 1'b1 ;
        16'd668 : reg_write_668 = 1'b1 ;
        16'd669 : reg_write_669 = 1'b1 ;
        16'd670 : reg_write_670 = 1'b1 ;
        16'd671 : reg_write_671 = 1'b1 ;
        16'd672 : reg_write_672 = 1'b1 ;
        16'd673 : reg_write_673 = 1'b1 ;
        16'd674 : reg_write_674 = 1'b1 ;
        16'd675 : reg_write_675 = 1'b1 ;
        16'd676 : reg_write_676 = 1'b1 ;
        16'd677 : reg_write_677 = 1'b1 ;
        16'd678 : reg_write_678 = 1'b1 ;
        16'd679 : reg_write_679 = 1'b1 ;
        16'd680 : reg_write_680 = 1'b1 ;
        16'd681 : reg_write_681 = 1'b1 ;
        16'd682 : reg_write_682 = 1'b1 ;
        16'd683 : reg_write_683 = 1'b1 ;
        16'd684 : reg_write_684 = 1'b1 ;
        16'd685 : reg_write_685 = 1'b1 ;
        16'd686 : reg_write_686 = 1'b1 ;
        16'd687 : reg_write_687 = 1'b1 ;
        16'd688 : reg_write_688 = 1'b1 ;
        16'd689 : reg_write_689 = 1'b1 ;
        16'd690 : reg_write_690 = 1'b1 ;
        16'd691 : reg_write_691 = 1'b1 ;
        16'd692 : reg_write_692 = 1'b1 ;
        16'd693 : reg_write_693 = 1'b1 ;
        16'd694 : reg_write_694 = 1'b1 ;
        16'd695 : reg_write_695 = 1'b1 ;
        16'd696 : reg_write_696 = 1'b1 ;
        16'd697 : reg_write_697 = 1'b1 ;
        16'd698 : reg_write_698 = 1'b1 ;
        16'd699 : reg_write_699 = 1'b1 ;
        16'd700 : reg_write_700 = 1'b1 ;
        16'd701 : reg_write_701 = 1'b1 ;
        16'd702 : reg_write_702 = 1'b1 ;
        16'd703 : reg_write_703 = 1'b1 ;
        16'd704 : reg_write_704 = 1'b1 ;
        16'd705 : reg_write_705 = 1'b1 ;
        16'd706 : reg_write_706 = 1'b1 ;
        16'd707 : reg_write_707 = 1'b1 ;
        16'd708 : reg_write_708 = 1'b1 ;
        16'd709 : reg_write_709 = 1'b1 ;
        16'd710 : reg_write_710 = 1'b1 ;
        16'd711 : reg_write_711 = 1'b1 ;
        16'd712 : reg_write_712 = 1'b1 ;
        16'd713 : reg_write_713 = 1'b1 ;
        16'd714 : reg_write_714 = 1'b1 ;
        16'd715 : reg_write_715 = 1'b1 ;
        16'd716 : reg_write_716 = 1'b1 ;
        16'd717 : reg_write_717 = 1'b1 ;
        16'd718 : reg_write_718 = 1'b1 ;
        16'd719 : reg_write_719 = 1'b1 ;
        16'd720 : reg_write_720 = 1'b1 ;
        16'd721 : reg_write_721 = 1'b1 ;
        16'd722 : reg_write_722 = 1'b1 ;
        16'd723 : reg_write_723 = 1'b1 ;
        16'd724 : reg_write_724 = 1'b1 ;
        16'd725 : reg_write_725 = 1'b1 ;
        16'd726 : reg_write_726 = 1'b1 ;
        16'd727 : reg_write_727 = 1'b1 ;
        16'd728 : reg_write_728 = 1'b1 ;
        16'd729 : reg_write_729 = 1'b1 ;
        16'd730 : reg_write_730 = 1'b1 ;
        16'd731 : reg_write_731 = 1'b1 ;
        16'd732 : reg_write_732 = 1'b1 ;
        16'd733 : reg_write_733 = 1'b1 ;
        16'd734 : reg_write_734 = 1'b1 ;
        16'd735 : reg_write_735 = 1'b1 ;
        16'd736 : reg_write_736 = 1'b1 ;
        16'd737 : reg_write_737 = 1'b1 ;
        16'd738 : reg_write_738 = 1'b1 ;
        16'd739 : reg_write_739 = 1'b1 ;
        16'd740 : reg_write_740 = 1'b1 ;
        16'd741 : reg_write_741 = 1'b1 ;
        16'd742 : reg_write_742 = 1'b1 ;
        16'd743 : reg_write_743 = 1'b1 ;
        16'd744 : reg_write_744 = 1'b1 ;
        16'd745 : reg_write_745 = 1'b1 ;
        16'd746 : reg_write_746 = 1'b1 ;
        16'd747 : reg_write_747 = 1'b1 ;
        16'd748 : reg_write_748 = 1'b1 ;
        16'd749 : reg_write_749 = 1'b1 ;
        16'd750 : reg_write_750 = 1'b1 ;
        16'd751 : reg_write_751 = 1'b1 ;
        16'd752 : reg_write_752 = 1'b1 ;
        16'd753 : reg_write_753 = 1'b1 ;
        16'd754 : reg_write_754 = 1'b1 ;
        16'd755 : reg_write_755 = 1'b1 ;
        16'd756 : reg_write_756 = 1'b1 ;
        16'd757 : reg_write_757 = 1'b1 ;
        16'd758 : reg_write_758 = 1'b1 ;
        16'd759 : reg_write_759 = 1'b1 ;
        16'd760 : reg_write_760 = 1'b1 ;
        16'd761 : reg_write_761 = 1'b1 ;
        16'd762 : reg_write_762 = 1'b1 ;
        16'd763 : reg_write_763 = 1'b1 ;
        16'd764 : reg_write_764 = 1'b1 ;
        16'd765 : reg_write_765 = 1'b1 ;
        16'd766 : reg_write_766 = 1'b1 ;
        16'd767 : reg_write_767 = 1'b1 ;
        16'd768 : reg_write_768 = 1'b1 ;
        16'd769 : reg_write_769 = 1'b1 ;
        16'd770 : reg_write_770 = 1'b1 ;
        16'd771 : reg_write_771 = 1'b1 ;
        16'd772 : reg_write_772 = 1'b1 ;
        16'd773 : reg_write_773 = 1'b1 ;
        16'd774 : reg_write_774 = 1'b1 ;
        16'd775 : reg_write_775 = 1'b1 ;
        16'd776 : reg_write_776 = 1'b1 ;
        16'd777 : reg_write_777 = 1'b1 ;
        16'd778 : reg_write_778 = 1'b1 ;
        16'd779 : reg_write_779 = 1'b1 ;
        16'd780 : reg_write_780 = 1'b1 ;
        16'd781 : reg_write_781 = 1'b1 ;
        16'd782 : reg_write_782 = 1'b1 ;
        16'd783 : reg_write_783 = 1'b1 ;
        16'd784 : reg_write_784 = 1'b1 ;
        16'd785 : reg_write_785 = 1'b1 ;
        16'd786 : reg_write_786 = 1'b1 ;
        16'd787 : reg_write_787 = 1'b1 ;
        16'd788 : reg_write_788 = 1'b1 ;
        16'd789 : reg_write_789 = 1'b1 ;
        16'd790 : reg_write_790 = 1'b1 ;
        16'd791 : reg_write_791 = 1'b1 ;
        16'd792 : reg_write_792 = 1'b1 ;
        16'd793 : reg_write_793 = 1'b1 ;
        16'd794 : reg_write_794 = 1'b1 ;
        16'd795 : reg_write_795 = 1'b1 ;
        16'd796 : reg_write_796 = 1'b1 ;
        16'd797 : reg_write_797 = 1'b1 ;
        16'd798 : reg_write_798 = 1'b1 ;
        16'd799 : reg_write_799 = 1'b1 ;
        16'd800 : reg_write_800 = 1'b1 ;
        16'd801 : reg_write_801 = 1'b1 ;
        16'd802 : reg_write_802 = 1'b1 ;
        16'd803 : reg_write_803 = 1'b1 ;
        16'd804 : reg_write_804 = 1'b1 ;
        16'd805 : reg_write_805 = 1'b1 ;
        16'd806 : reg_write_806 = 1'b1 ;
        16'd807 : reg_write_807 = 1'b1 ;
        16'd808 : reg_write_808 = 1'b1 ;
        16'd809 : reg_write_809 = 1'b1 ;
        16'd810 : reg_write_810 = 1'b1 ;
        16'd811 : reg_write_811 = 1'b1 ;
        16'd812 : reg_write_812 = 1'b1 ;
        16'd813 : reg_write_813 = 1'b1 ;
        16'd814 : reg_write_814 = 1'b1 ;
        16'd815 : reg_write_815 = 1'b1 ;
        16'd816 : reg_write_816 = 1'b1 ;
        16'd817 : reg_write_817 = 1'b1 ;
        16'd818 : reg_write_818 = 1'b1 ;
        16'd819 : reg_write_819 = 1'b1 ;
        16'd820 : reg_write_820 = 1'b1 ;
        16'd821 : reg_write_821 = 1'b1 ;
        16'd822 : reg_write_822 = 1'b1 ;
        16'd823 : reg_write_823 = 1'b1 ;
        16'd824 : reg_write_824 = 1'b1 ;
        16'd825 : reg_write_825 = 1'b1 ;
        16'd826 : reg_write_826 = 1'b1 ;
        16'd827 : reg_write_827 = 1'b1 ;
        16'd828 : reg_write_828 = 1'b1 ;
        16'd829 : reg_write_829 = 1'b1 ;
        16'd830 : reg_write_830 = 1'b1 ;
        16'd831 : reg_write_831 = 1'b1 ;
        16'd832 : reg_write_832 = 1'b1 ;
        16'd833 : reg_write_833 = 1'b1 ;
        16'd834 : reg_write_834 = 1'b1 ;
        16'd835 : reg_write_835 = 1'b1 ;
        16'd836 : reg_write_836 = 1'b1 ;
        16'd837 : reg_write_837 = 1'b1 ;
        16'd838 : reg_write_838 = 1'b1 ;
        16'd839 : reg_write_839 = 1'b1 ;
        16'd840 : reg_write_840 = 1'b1 ;
        16'd841 : reg_write_841 = 1'b1 ;
        16'd842 : reg_write_842 = 1'b1 ;
        16'd843 : reg_write_843 = 1'b1 ;
        16'd844 : reg_write_844 = 1'b1 ;
        16'd845 : reg_write_845 = 1'b1 ;
        16'd846 : reg_write_846 = 1'b1 ;
        16'd847 : reg_write_847 = 1'b1 ;
        16'd848 : reg_write_848 = 1'b1 ;
        16'd849 : reg_write_849 = 1'b1 ;
        16'd850 : reg_write_850 = 1'b1 ;
        16'd851 : reg_write_851 = 1'b1 ;
        16'd852 : reg_write_852 = 1'b1 ;
        16'd853 : reg_write_853 = 1'b1 ;
        16'd854 : reg_write_854 = 1'b1 ;
        16'd855 : reg_write_855 = 1'b1 ;
        16'd856 : reg_write_856 = 1'b1 ;
        16'd857 : reg_write_857 = 1'b1 ;
        16'd858 : reg_write_858 = 1'b1 ;
        16'd859 : reg_write_859 = 1'b1 ;
        16'd860 : reg_write_860 = 1'b1 ;
        16'd861 : reg_write_861 = 1'b1 ;
        16'd862 : reg_write_862 = 1'b1 ;
        16'd863 : reg_write_863 = 1'b1 ;
        16'd864 : reg_write_864 = 1'b1 ;
        16'd865 : reg_write_865 = 1'b1 ;
        16'd866 : reg_write_866 = 1'b1 ;
        16'd867 : reg_write_867 = 1'b1 ;
        16'd868 : reg_write_868 = 1'b1 ;
        16'd869 : reg_write_869 = 1'b1 ;
        16'd870 : reg_write_870 = 1'b1 ;
        16'd871 : reg_write_871 = 1'b1 ;
        16'd872 : reg_write_872 = 1'b1 ;
        16'd873 : reg_write_873 = 1'b1 ;
        16'd874 : reg_write_874 = 1'b1 ;
        16'd875 : reg_write_875 = 1'b1 ;
        16'd876 : reg_write_876 = 1'b1 ;
        16'd877 : reg_write_877 = 1'b1 ;
        16'd878 : reg_write_878 = 1'b1 ;
        16'd879 : reg_write_879 = 1'b1 ;
        16'd880 : reg_write_880 = 1'b1 ;
        16'd881 : reg_write_881 = 1'b1 ;
        16'd882 : reg_write_882 = 1'b1 ;
        16'd883 : reg_write_883 = 1'b1 ;
        16'd884 : reg_write_884 = 1'b1 ;
        16'd885 : reg_write_885 = 1'b1 ;
        16'd886 : reg_write_886 = 1'b1 ;
        16'd887 : reg_write_887 = 1'b1 ;
        16'd888 : reg_write_888 = 1'b1 ;
        16'd889 : reg_write_889 = 1'b1 ;
        16'd890 : reg_write_890 = 1'b1 ;
        16'd891 : reg_write_891 = 1'b1 ;
        16'd892 : reg_write_892 = 1'b1 ;
        16'd893 : reg_write_893 = 1'b1 ;
        16'd894 : reg_write_894 = 1'b1 ;
        16'd895 : reg_write_895 = 1'b1 ;
        16'd896 : reg_write_896 = 1'b1 ;
        16'd897 : reg_write_897 = 1'b1 ;
        16'd898 : reg_write_898 = 1'b1 ;
        16'd899 : reg_write_899 = 1'b1 ;
        16'd900 : reg_write_900 = 1'b1 ;
        16'd901 : reg_write_901 = 1'b1 ;
        16'd902 : reg_write_902 = 1'b1 ;
        16'd903 : reg_write_903 = 1'b1 ;
        16'd904 : reg_write_904 = 1'b1 ;
        16'd905 : reg_write_905 = 1'b1 ;
        16'd906 : reg_write_906 = 1'b1 ;
        16'd907 : reg_write_907 = 1'b1 ;
        16'd908 : reg_write_908 = 1'b1 ;
        16'd909 : reg_write_909 = 1'b1 ;
        16'd910 : reg_write_910 = 1'b1 ;
        16'd911 : reg_write_911 = 1'b1 ;
        16'd912 : reg_write_912 = 1'b1 ;
        16'd913 : reg_write_913 = 1'b1 ;
        16'd914 : reg_write_914 = 1'b1 ;
        16'd915 : reg_write_915 = 1'b1 ;
        16'd916 : reg_write_916 = 1'b1 ;
        16'd917 : reg_write_917 = 1'b1 ;
        16'd918 : reg_write_918 = 1'b1 ;
        16'd919 : reg_write_919 = 1'b1 ;
        16'd920 : reg_write_920 = 1'b1 ;
        16'd921 : reg_write_921 = 1'b1 ;
        16'd922 : reg_write_922 = 1'b1 ;
        16'd923 : reg_write_923 = 1'b1 ;
        16'd924 : reg_write_924 = 1'b1 ;
        16'd925 : reg_write_925 = 1'b1 ;
        16'd926 : reg_write_926 = 1'b1 ;
        16'd927 : reg_write_927 = 1'b1 ;
        16'd928 : reg_write_928 = 1'b1 ;
        16'd929 : reg_write_929 = 1'b1 ;
        16'd930 : reg_write_930 = 1'b1 ;
        16'd931 : reg_write_931 = 1'b1 ;
        16'd932 : reg_write_932 = 1'b1 ;
        16'd933 : reg_write_933 = 1'b1 ;
        16'd934 : reg_write_934 = 1'b1 ;
        16'd935 : reg_write_935 = 1'b1 ;
        16'd936 : reg_write_936 = 1'b1 ;
        16'd937 : reg_write_937 = 1'b1 ;
        16'd938 : reg_write_938 = 1'b1 ;
        16'd939 : reg_write_939 = 1'b1 ;
        16'd940 : reg_write_940 = 1'b1 ;
        16'd941 : reg_write_941 = 1'b1 ;
        16'd942 : reg_write_942 = 1'b1 ;
        16'd943 : reg_write_943 = 1'b1 ;
        16'd944 : reg_write_944 = 1'b1 ;
        16'd945 : reg_write_945 = 1'b1 ;
        16'd946 : reg_write_946 = 1'b1 ;
        16'd947 : reg_write_947 = 1'b1 ;
        16'd948 : reg_write_948 = 1'b1 ;
        16'd949 : reg_write_949 = 1'b1 ;
        16'd950 : reg_write_950 = 1'b1 ;
        16'd951 : reg_write_951 = 1'b1 ;
        16'd952 : reg_write_952 = 1'b1 ;
        16'd953 : reg_write_953 = 1'b1 ;
        16'd954 : reg_write_954 = 1'b1 ;
        16'd955 : reg_write_955 = 1'b1 ;
        16'd956 : reg_write_956 = 1'b1 ;
        16'd957 : reg_write_957 = 1'b1 ;
        16'd958 : reg_write_958 = 1'b1 ;
        16'd959 : reg_write_959 = 1'b1 ;
        16'd960 : reg_write_960 = 1'b1 ;
        16'd961 : reg_write_961 = 1'b1 ;
        16'd962 : reg_write_962 = 1'b1 ;
        16'd963 : reg_write_963 = 1'b1 ;
        16'd964 : reg_write_964 = 1'b1 ;
        16'd965 : reg_write_965 = 1'b1 ;
        16'd966 : reg_write_966 = 1'b1 ;
        16'd967 : reg_write_967 = 1'b1 ;
        16'd968 : reg_write_968 = 1'b1 ;
        16'd969 : reg_write_969 = 1'b1 ;
        16'd970 : reg_write_970 = 1'b1 ;
        16'd971 : reg_write_971 = 1'b1 ;
        16'd972 : reg_write_972 = 1'b1 ;
        16'd973 : reg_write_973 = 1'b1 ;
        16'd974 : reg_write_974 = 1'b1 ;
        16'd975 : reg_write_975 = 1'b1 ;
        16'd976 : reg_write_976 = 1'b1 ;
        16'd977 : reg_write_977 = 1'b1 ;
        16'd978 : reg_write_978 = 1'b1 ;
        16'd979 : reg_write_979 = 1'b1 ;
        16'd980 : reg_write_980 = 1'b1 ;
        16'd981 : reg_write_981 = 1'b1 ;
        16'd982 : reg_write_982 = 1'b1 ;
        16'd983 : reg_write_983 = 1'b1 ;
        16'd984 : reg_write_984 = 1'b1 ;
        16'd985 : reg_write_985 = 1'b1 ;
        16'd986 : reg_write_986 = 1'b1 ;
        16'd987 : reg_write_987 = 1'b1 ;
        16'd988 : reg_write_988 = 1'b1 ;
        16'd989 : reg_write_989 = 1'b1 ;
        16'd990 : reg_write_990 = 1'b1 ;
        16'd991 : reg_write_991 = 1'b1 ;
        16'd992 : reg_write_992 = 1'b1 ;
        16'd993 : reg_write_993 = 1'b1 ;
        16'd994 : reg_write_994 = 1'b1 ;
        16'd995 : reg_write_995 = 1'b1 ;
        16'd996 : reg_write_996 = 1'b1 ;
        16'd997 : reg_write_997 = 1'b1 ;
        16'd998 : reg_write_998 = 1'b1 ;
        16'd999 : reg_write_999 = 1'b1 ;
        16'd1000 : reg_write_1000 = 1'b1 ;
			endcase 
			end
			else begin
        reg_write_1 = 1'b0 ;
        reg_write_2 = 1'b0 ;
        reg_write_3 = 1'b0 ;
        reg_write_4 = 1'b0 ;
        reg_write_5 = 1'b0 ;
        reg_write_6 = 1'b0 ;
        reg_write_7 = 1'b0 ;
        reg_write_8 = 1'b0 ;
        reg_write_9 = 1'b0 ;
        reg_write_10 = 1'b0 ;
        reg_write_11 = 1'b0 ;
        reg_write_12 = 1'b0 ;
        reg_write_13 = 1'b0 ;
        reg_write_14 = 1'b0 ;
        reg_write_15 = 1'b0 ;
        reg_write_16 = 1'b0 ;
        reg_write_17 = 1'b0 ;
        reg_write_18 = 1'b0 ;
        reg_write_19 = 1'b0 ;
        reg_write_20 = 1'b0 ;
        reg_write_21 = 1'b0 ;
        reg_write_22 = 1'b0 ;
        reg_write_23 = 1'b0 ;
        reg_write_24 = 1'b0 ;
        reg_write_25 = 1'b0 ;
        reg_write_26 = 1'b0 ;
        reg_write_27 = 1'b0 ;
        reg_write_28 = 1'b0 ;
        reg_write_29 = 1'b0 ;
        reg_write_30 = 1'b0 ;
        reg_write_31 = 1'b0 ;
        reg_write_32 = 1'b0 ;
        reg_write_33 = 1'b0 ;
        reg_write_34 = 1'b0 ;
        reg_write_35 = 1'b0 ;
        reg_write_36 = 1'b0 ;
        reg_write_37 = 1'b0 ;
        reg_write_38 = 1'b0 ;
        reg_write_39 = 1'b0 ;
        reg_write_40 = 1'b0 ;
        reg_write_41 = 1'b0 ;
        reg_write_42 = 1'b0 ;
        reg_write_43 = 1'b0 ;
        reg_write_44 = 1'b0 ;
        reg_write_45 = 1'b0 ;
        reg_write_46 = 1'b0 ;
        reg_write_47 = 1'b0 ;
        reg_write_48 = 1'b0 ;
        reg_write_49 = 1'b0 ;
        reg_write_50 = 1'b0 ;
        reg_write_51 = 1'b0 ;
        reg_write_52 = 1'b0 ;
        reg_write_53 = 1'b0 ;
        reg_write_54 = 1'b0 ;
        reg_write_55 = 1'b0 ;
        reg_write_56 = 1'b0 ;
        reg_write_57 = 1'b0 ;
        reg_write_58 = 1'b0 ;
        reg_write_59 = 1'b0 ;
        reg_write_60 = 1'b0 ;
        reg_write_61 = 1'b0 ;
        reg_write_62 = 1'b0 ;
        reg_write_63 = 1'b0 ;
        reg_write_64 = 1'b0 ;
        reg_write_65 = 1'b0 ;
        reg_write_66 = 1'b0 ;
        reg_write_67 = 1'b0 ;
        reg_write_68 = 1'b0 ;
        reg_write_69 = 1'b0 ;
        reg_write_70 = 1'b0 ;
        reg_write_71 = 1'b0 ;
        reg_write_72 = 1'b0 ;
        reg_write_73 = 1'b0 ;
        reg_write_74 = 1'b0 ;
        reg_write_75 = 1'b0 ;
        reg_write_76 = 1'b0 ;
        reg_write_77 = 1'b0 ;
        reg_write_78 = 1'b0 ;
        reg_write_79 = 1'b0 ;
        reg_write_80 = 1'b0 ;
        reg_write_81 = 1'b0 ;
        reg_write_82 = 1'b0 ;
        reg_write_83 = 1'b0 ;
        reg_write_84 = 1'b0 ;
        reg_write_85 = 1'b0 ;
        reg_write_86 = 1'b0 ;
        reg_write_87 = 1'b0 ;
        reg_write_88 = 1'b0 ;
        reg_write_89 = 1'b0 ;
        reg_write_90 = 1'b0 ;
        reg_write_91 = 1'b0 ;
        reg_write_92 = 1'b0 ;
        reg_write_93 = 1'b0 ;
        reg_write_94 = 1'b0 ;
        reg_write_95 = 1'b0 ;
        reg_write_96 = 1'b0 ;
        reg_write_97 = 1'b0 ;
        reg_write_98 = 1'b0 ;
        reg_write_99 = 1'b0 ;
        reg_write_100 = 1'b0 ;
        reg_write_101 = 1'b0 ;
        reg_write_102 = 1'b0 ;
        reg_write_103 = 1'b0 ;
        reg_write_104 = 1'b0 ;
        reg_write_105 = 1'b0 ;
        reg_write_106 = 1'b0 ;
        reg_write_107 = 1'b0 ;
        reg_write_108 = 1'b0 ;
        reg_write_109 = 1'b0 ;
        reg_write_110 = 1'b0 ;
        reg_write_111 = 1'b0 ;
        reg_write_112 = 1'b0 ;
        reg_write_113 = 1'b0 ;
        reg_write_114 = 1'b0 ;
        reg_write_115 = 1'b0 ;
        reg_write_116 = 1'b0 ;
        reg_write_117 = 1'b0 ;
        reg_write_118 = 1'b0 ;
        reg_write_119 = 1'b0 ;
        reg_write_120 = 1'b0 ;
        reg_write_121 = 1'b0 ;
        reg_write_122 = 1'b0 ;
        reg_write_123 = 1'b0 ;
        reg_write_124 = 1'b0 ;
        reg_write_125 = 1'b0 ;
        reg_write_126 = 1'b0 ;
        reg_write_127 = 1'b0 ;
        reg_write_128 = 1'b0 ;
        reg_write_129 = 1'b0 ;
        reg_write_130 = 1'b0 ;
        reg_write_131 = 1'b0 ;
        reg_write_132 = 1'b0 ;
        reg_write_133 = 1'b0 ;
        reg_write_134 = 1'b0 ;
        reg_write_135 = 1'b0 ;
        reg_write_136 = 1'b0 ;
        reg_write_137 = 1'b0 ;
        reg_write_138 = 1'b0 ;
        reg_write_139 = 1'b0 ;
        reg_write_140 = 1'b0 ;
        reg_write_141 = 1'b0 ;
        reg_write_142 = 1'b0 ;
        reg_write_143 = 1'b0 ;
        reg_write_144 = 1'b0 ;
        reg_write_145 = 1'b0 ;
        reg_write_146 = 1'b0 ;
        reg_write_147 = 1'b0 ;
        reg_write_148 = 1'b0 ;
        reg_write_149 = 1'b0 ;
        reg_write_150 = 1'b0 ;
        reg_write_151 = 1'b0 ;
        reg_write_152 = 1'b0 ;
        reg_write_153 = 1'b0 ;
        reg_write_154 = 1'b0 ;
        reg_write_155 = 1'b0 ;
        reg_write_156 = 1'b0 ;
        reg_write_157 = 1'b0 ;
        reg_write_158 = 1'b0 ;
        reg_write_159 = 1'b0 ;
        reg_write_160 = 1'b0 ;
        reg_write_161 = 1'b0 ;
        reg_write_162 = 1'b0 ;
        reg_write_163 = 1'b0 ;
        reg_write_164 = 1'b0 ;
        reg_write_165 = 1'b0 ;
        reg_write_166 = 1'b0 ;
        reg_write_167 = 1'b0 ;
        reg_write_168 = 1'b0 ;
        reg_write_169 = 1'b0 ;
        reg_write_170 = 1'b0 ;
        reg_write_171 = 1'b0 ;
        reg_write_172 = 1'b0 ;
        reg_write_173 = 1'b0 ;
        reg_write_174 = 1'b0 ;
        reg_write_175 = 1'b0 ;
        reg_write_176 = 1'b0 ;
        reg_write_177 = 1'b0 ;
        reg_write_178 = 1'b0 ;
        reg_write_179 = 1'b0 ;
        reg_write_180 = 1'b0 ;
        reg_write_181 = 1'b0 ;
        reg_write_182 = 1'b0 ;
        reg_write_183 = 1'b0 ;
        reg_write_184 = 1'b0 ;
        reg_write_185 = 1'b0 ;
        reg_write_186 = 1'b0 ;
        reg_write_187 = 1'b0 ;
        reg_write_188 = 1'b0 ;
        reg_write_189 = 1'b0 ;
        reg_write_190 = 1'b0 ;
        reg_write_191 = 1'b0 ;
        reg_write_192 = 1'b0 ;
        reg_write_193 = 1'b0 ;
        reg_write_194 = 1'b0 ;
        reg_write_195 = 1'b0 ;
        reg_write_196 = 1'b0 ;
        reg_write_197 = 1'b0 ;
        reg_write_198 = 1'b0 ;
        reg_write_199 = 1'b0 ;
        reg_write_200 = 1'b0 ;
        reg_write_201 = 1'b0 ;
        reg_write_202 = 1'b0 ;
        reg_write_203 = 1'b0 ;
        reg_write_204 = 1'b0 ;
        reg_write_205 = 1'b0 ;
        reg_write_206 = 1'b0 ;
        reg_write_207 = 1'b0 ;
        reg_write_208 = 1'b0 ;
        reg_write_209 = 1'b0 ;
        reg_write_210 = 1'b0 ;
        reg_write_211 = 1'b0 ;
        reg_write_212 = 1'b0 ;
        reg_write_213 = 1'b0 ;
        reg_write_214 = 1'b0 ;
        reg_write_215 = 1'b0 ;
        reg_write_216 = 1'b0 ;
        reg_write_217 = 1'b0 ;
        reg_write_218 = 1'b0 ;
        reg_write_219 = 1'b0 ;
        reg_write_220 = 1'b0 ;
        reg_write_221 = 1'b0 ;
        reg_write_222 = 1'b0 ;
        reg_write_223 = 1'b0 ;
        reg_write_224 = 1'b0 ;
        reg_write_225 = 1'b0 ;
        reg_write_226 = 1'b0 ;
        reg_write_227 = 1'b0 ;
        reg_write_228 = 1'b0 ;
        reg_write_229 = 1'b0 ;
        reg_write_230 = 1'b0 ;
        reg_write_231 = 1'b0 ;
        reg_write_232 = 1'b0 ;
        reg_write_233 = 1'b0 ;
        reg_write_234 = 1'b0 ;
        reg_write_235 = 1'b0 ;
        reg_write_236 = 1'b0 ;
        reg_write_237 = 1'b0 ;
        reg_write_238 = 1'b0 ;
        reg_write_239 = 1'b0 ;
        reg_write_240 = 1'b0 ;
        reg_write_241 = 1'b0 ;
        reg_write_242 = 1'b0 ;
        reg_write_243 = 1'b0 ;
        reg_write_244 = 1'b0 ;
        reg_write_245 = 1'b0 ;
        reg_write_246 = 1'b0 ;
        reg_write_247 = 1'b0 ;
        reg_write_248 = 1'b0 ;
        reg_write_249 = 1'b0 ;
        reg_write_250 = 1'b0 ;
        reg_write_251 = 1'b0 ;
        reg_write_252 = 1'b0 ;
        reg_write_253 = 1'b0 ;
        reg_write_254 = 1'b0 ;
        reg_write_255 = 1'b0 ;
        reg_write_256 = 1'b0 ;
        reg_write_257 = 1'b0 ;
        reg_write_258 = 1'b0 ;
        reg_write_259 = 1'b0 ;
        reg_write_260 = 1'b0 ;
        reg_write_261 = 1'b0 ;
        reg_write_262 = 1'b0 ;
        reg_write_263 = 1'b0 ;
        reg_write_264 = 1'b0 ;
        reg_write_265 = 1'b0 ;
        reg_write_266 = 1'b0 ;
        reg_write_267 = 1'b0 ;
        reg_write_268 = 1'b0 ;
        reg_write_269 = 1'b0 ;
        reg_write_270 = 1'b0 ;
        reg_write_271 = 1'b0 ;
        reg_write_272 = 1'b0 ;
        reg_write_273 = 1'b0 ;
        reg_write_274 = 1'b0 ;
        reg_write_275 = 1'b0 ;
        reg_write_276 = 1'b0 ;
        reg_write_277 = 1'b0 ;
        reg_write_278 = 1'b0 ;
        reg_write_279 = 1'b0 ;
        reg_write_280 = 1'b0 ;
        reg_write_281 = 1'b0 ;
        reg_write_282 = 1'b0 ;
        reg_write_283 = 1'b0 ;
        reg_write_284 = 1'b0 ;
        reg_write_285 = 1'b0 ;
        reg_write_286 = 1'b0 ;
        reg_write_287 = 1'b0 ;
        reg_write_288 = 1'b0 ;
        reg_write_289 = 1'b0 ;
        reg_write_290 = 1'b0 ;
        reg_write_291 = 1'b0 ;
        reg_write_292 = 1'b0 ;
        reg_write_293 = 1'b0 ;
        reg_write_294 = 1'b0 ;
        reg_write_295 = 1'b0 ;
        reg_write_296 = 1'b0 ;
        reg_write_297 = 1'b0 ;
        reg_write_298 = 1'b0 ;
        reg_write_299 = 1'b0 ;
        reg_write_300 = 1'b0 ;
        reg_write_301 = 1'b0 ;
        reg_write_302 = 1'b0 ;
        reg_write_303 = 1'b0 ;
        reg_write_304 = 1'b0 ;
        reg_write_305 = 1'b0 ;
        reg_write_306 = 1'b0 ;
        reg_write_307 = 1'b0 ;
        reg_write_308 = 1'b0 ;
        reg_write_309 = 1'b0 ;
        reg_write_310 = 1'b0 ;
        reg_write_311 = 1'b0 ;
        reg_write_312 = 1'b0 ;
        reg_write_313 = 1'b0 ;
        reg_write_314 = 1'b0 ;
        reg_write_315 = 1'b0 ;
        reg_write_316 = 1'b0 ;
        reg_write_317 = 1'b0 ;
        reg_write_318 = 1'b0 ;
        reg_write_319 = 1'b0 ;
        reg_write_320 = 1'b0 ;
        reg_write_321 = 1'b0 ;
        reg_write_322 = 1'b0 ;
        reg_write_323 = 1'b0 ;
        reg_write_324 = 1'b0 ;
        reg_write_325 = 1'b0 ;
        reg_write_326 = 1'b0 ;
        reg_write_327 = 1'b0 ;
        reg_write_328 = 1'b0 ;
        reg_write_329 = 1'b0 ;
        reg_write_330 = 1'b0 ;
        reg_write_331 = 1'b0 ;
        reg_write_332 = 1'b0 ;
        reg_write_333 = 1'b0 ;
        reg_write_334 = 1'b0 ;
        reg_write_335 = 1'b0 ;
        reg_write_336 = 1'b0 ;
        reg_write_337 = 1'b0 ;
        reg_write_338 = 1'b0 ;
        reg_write_339 = 1'b0 ;
        reg_write_340 = 1'b0 ;
        reg_write_341 = 1'b0 ;
        reg_write_342 = 1'b0 ;
        reg_write_343 = 1'b0 ;
        reg_write_344 = 1'b0 ;
        reg_write_345 = 1'b0 ;
        reg_write_346 = 1'b0 ;
        reg_write_347 = 1'b0 ;
        reg_write_348 = 1'b0 ;
        reg_write_349 = 1'b0 ;
        reg_write_350 = 1'b0 ;
        reg_write_351 = 1'b0 ;
        reg_write_352 = 1'b0 ;
        reg_write_353 = 1'b0 ;
        reg_write_354 = 1'b0 ;
        reg_write_355 = 1'b0 ;
        reg_write_356 = 1'b0 ;
        reg_write_357 = 1'b0 ;
        reg_write_358 = 1'b0 ;
        reg_write_359 = 1'b0 ;
        reg_write_360 = 1'b0 ;
        reg_write_361 = 1'b0 ;
        reg_write_362 = 1'b0 ;
        reg_write_363 = 1'b0 ;
        reg_write_364 = 1'b0 ;
        reg_write_365 = 1'b0 ;
        reg_write_366 = 1'b0 ;
        reg_write_367 = 1'b0 ;
        reg_write_368 = 1'b0 ;
        reg_write_369 = 1'b0 ;
        reg_write_370 = 1'b0 ;
        reg_write_371 = 1'b0 ;
        reg_write_372 = 1'b0 ;
        reg_write_373 = 1'b0 ;
        reg_write_374 = 1'b0 ;
        reg_write_375 = 1'b0 ;
        reg_write_376 = 1'b0 ;
        reg_write_377 = 1'b0 ;
        reg_write_378 = 1'b0 ;
        reg_write_379 = 1'b0 ;
        reg_write_380 = 1'b0 ;
        reg_write_381 = 1'b0 ;
        reg_write_382 = 1'b0 ;
        reg_write_383 = 1'b0 ;
        reg_write_384 = 1'b0 ;
        reg_write_385 = 1'b0 ;
        reg_write_386 = 1'b0 ;
        reg_write_387 = 1'b0 ;
        reg_write_388 = 1'b0 ;
        reg_write_389 = 1'b0 ;
        reg_write_390 = 1'b0 ;
        reg_write_391 = 1'b0 ;
        reg_write_392 = 1'b0 ;
        reg_write_393 = 1'b0 ;
        reg_write_394 = 1'b0 ;
        reg_write_395 = 1'b0 ;
        reg_write_396 = 1'b0 ;
        reg_write_397 = 1'b0 ;
        reg_write_398 = 1'b0 ;
        reg_write_399 = 1'b0 ;
        reg_write_400 = 1'b0 ;
        reg_write_401 = 1'b0 ;
        reg_write_402 = 1'b0 ;
        reg_write_403 = 1'b0 ;
        reg_write_404 = 1'b0 ;
        reg_write_405 = 1'b0 ;
        reg_write_406 = 1'b0 ;
        reg_write_407 = 1'b0 ;
        reg_write_408 = 1'b0 ;
        reg_write_409 = 1'b0 ;
        reg_write_410 = 1'b0 ;
        reg_write_411 = 1'b0 ;
        reg_write_412 = 1'b0 ;
        reg_write_413 = 1'b0 ;
        reg_write_414 = 1'b0 ;
        reg_write_415 = 1'b0 ;
        reg_write_416 = 1'b0 ;
        reg_write_417 = 1'b0 ;
        reg_write_418 = 1'b0 ;
        reg_write_419 = 1'b0 ;
        reg_write_420 = 1'b0 ;
        reg_write_421 = 1'b0 ;
        reg_write_422 = 1'b0 ;
        reg_write_423 = 1'b0 ;
        reg_write_424 = 1'b0 ;
        reg_write_425 = 1'b0 ;
        reg_write_426 = 1'b0 ;
        reg_write_427 = 1'b0 ;
        reg_write_428 = 1'b0 ;
        reg_write_429 = 1'b0 ;
        reg_write_430 = 1'b0 ;
        reg_write_431 = 1'b0 ;
        reg_write_432 = 1'b0 ;
        reg_write_433 = 1'b0 ;
        reg_write_434 = 1'b0 ;
        reg_write_435 = 1'b0 ;
        reg_write_436 = 1'b0 ;
        reg_write_437 = 1'b0 ;
        reg_write_438 = 1'b0 ;
        reg_write_439 = 1'b0 ;
        reg_write_440 = 1'b0 ;
        reg_write_441 = 1'b0 ;
        reg_write_442 = 1'b0 ;
        reg_write_443 = 1'b0 ;
        reg_write_444 = 1'b0 ;
        reg_write_445 = 1'b0 ;
        reg_write_446 = 1'b0 ;
        reg_write_447 = 1'b0 ;
        reg_write_448 = 1'b0 ;
        reg_write_449 = 1'b0 ;
        reg_write_450 = 1'b0 ;
        reg_write_451 = 1'b0 ;
        reg_write_452 = 1'b0 ;
        reg_write_453 = 1'b0 ;
        reg_write_454 = 1'b0 ;
        reg_write_455 = 1'b0 ;
        reg_write_456 = 1'b0 ;
        reg_write_457 = 1'b0 ;
        reg_write_458 = 1'b0 ;
        reg_write_459 = 1'b0 ;
        reg_write_460 = 1'b0 ;
        reg_write_461 = 1'b0 ;
        reg_write_462 = 1'b0 ;
        reg_write_463 = 1'b0 ;
        reg_write_464 = 1'b0 ;
        reg_write_465 = 1'b0 ;
        reg_write_466 = 1'b0 ;
        reg_write_467 = 1'b0 ;
        reg_write_468 = 1'b0 ;
        reg_write_469 = 1'b0 ;
        reg_write_470 = 1'b0 ;
        reg_write_471 = 1'b0 ;
        reg_write_472 = 1'b0 ;
        reg_write_473 = 1'b0 ;
        reg_write_474 = 1'b0 ;
        reg_write_475 = 1'b0 ;
        reg_write_476 = 1'b0 ;
        reg_write_477 = 1'b0 ;
        reg_write_478 = 1'b0 ;
        reg_write_479 = 1'b0 ;
        reg_write_480 = 1'b0 ;
        reg_write_481 = 1'b0 ;
        reg_write_482 = 1'b0 ;
        reg_write_483 = 1'b0 ;
        reg_write_484 = 1'b0 ;
        reg_write_485 = 1'b0 ;
        reg_write_486 = 1'b0 ;
        reg_write_487 = 1'b0 ;
        reg_write_488 = 1'b0 ;
        reg_write_489 = 1'b0 ;
        reg_write_490 = 1'b0 ;
        reg_write_491 = 1'b0 ;
        reg_write_492 = 1'b0 ;
        reg_write_493 = 1'b0 ;
        reg_write_494 = 1'b0 ;
        reg_write_495 = 1'b0 ;
        reg_write_496 = 1'b0 ;
        reg_write_497 = 1'b0 ;
        reg_write_498 = 1'b0 ;
        reg_write_499 = 1'b0 ;
        reg_write_500 = 1'b0 ;
        reg_write_501 = 1'b0 ;
        reg_write_502 = 1'b0 ;
        reg_write_503 = 1'b0 ;
        reg_write_504 = 1'b0 ;
        reg_write_505 = 1'b0 ;
        reg_write_506 = 1'b0 ;
        reg_write_507 = 1'b0 ;
        reg_write_508 = 1'b0 ;
        reg_write_509 = 1'b0 ;
        reg_write_510 = 1'b0 ;
        reg_write_511 = 1'b0 ;
        reg_write_512 = 1'b0 ;
        reg_write_513 = 1'b0 ;
        reg_write_514 = 1'b0 ;
        reg_write_515 = 1'b0 ;
        reg_write_516 = 1'b0 ;
        reg_write_517 = 1'b0 ;
        reg_write_518 = 1'b0 ;
        reg_write_519 = 1'b0 ;
        reg_write_520 = 1'b0 ;
        reg_write_521 = 1'b0 ;
        reg_write_522 = 1'b0 ;
        reg_write_523 = 1'b0 ;
        reg_write_524 = 1'b0 ;
        reg_write_525 = 1'b0 ;
        reg_write_526 = 1'b0 ;
        reg_write_527 = 1'b0 ;
        reg_write_528 = 1'b0 ;
        reg_write_529 = 1'b0 ;
        reg_write_530 = 1'b0 ;
        reg_write_531 = 1'b0 ;
        reg_write_532 = 1'b0 ;
        reg_write_533 = 1'b0 ;
        reg_write_534 = 1'b0 ;
        reg_write_535 = 1'b0 ;
        reg_write_536 = 1'b0 ;
        reg_write_537 = 1'b0 ;
        reg_write_538 = 1'b0 ;
        reg_write_539 = 1'b0 ;
        reg_write_540 = 1'b0 ;
        reg_write_541 = 1'b0 ;
        reg_write_542 = 1'b0 ;
        reg_write_543 = 1'b0 ;
        reg_write_544 = 1'b0 ;
        reg_write_545 = 1'b0 ;
        reg_write_546 = 1'b0 ;
        reg_write_547 = 1'b0 ;
        reg_write_548 = 1'b0 ;
        reg_write_549 = 1'b0 ;
        reg_write_550 = 1'b0 ;
        reg_write_551 = 1'b0 ;
        reg_write_552 = 1'b0 ;
        reg_write_553 = 1'b0 ;
        reg_write_554 = 1'b0 ;
        reg_write_555 = 1'b0 ;
        reg_write_556 = 1'b0 ;
        reg_write_557 = 1'b0 ;
        reg_write_558 = 1'b0 ;
        reg_write_559 = 1'b0 ;
        reg_write_560 = 1'b0 ;
        reg_write_561 = 1'b0 ;
        reg_write_562 = 1'b0 ;
        reg_write_563 = 1'b0 ;
        reg_write_564 = 1'b0 ;
        reg_write_565 = 1'b0 ;
        reg_write_566 = 1'b0 ;
        reg_write_567 = 1'b0 ;
        reg_write_568 = 1'b0 ;
        reg_write_569 = 1'b0 ;
        reg_write_570 = 1'b0 ;
        reg_write_571 = 1'b0 ;
        reg_write_572 = 1'b0 ;
        reg_write_573 = 1'b0 ;
        reg_write_574 = 1'b0 ;
        reg_write_575 = 1'b0 ;
        reg_write_576 = 1'b0 ;
        reg_write_577 = 1'b0 ;
        reg_write_578 = 1'b0 ;
        reg_write_579 = 1'b0 ;
        reg_write_580 = 1'b0 ;
        reg_write_581 = 1'b0 ;
        reg_write_582 = 1'b0 ;
        reg_write_583 = 1'b0 ;
        reg_write_584 = 1'b0 ;
        reg_write_585 = 1'b0 ;
        reg_write_586 = 1'b0 ;
        reg_write_587 = 1'b0 ;
        reg_write_588 = 1'b0 ;
        reg_write_589 = 1'b0 ;
        reg_write_590 = 1'b0 ;
        reg_write_591 = 1'b0 ;
        reg_write_592 = 1'b0 ;
        reg_write_593 = 1'b0 ;
        reg_write_594 = 1'b0 ;
        reg_write_595 = 1'b0 ;
        reg_write_596 = 1'b0 ;
        reg_write_597 = 1'b0 ;
        reg_write_598 = 1'b0 ;
        reg_write_599 = 1'b0 ;
        reg_write_600 = 1'b0 ;
        reg_write_601 = 1'b0 ;
        reg_write_602 = 1'b0 ;
        reg_write_603 = 1'b0 ;
        reg_write_604 = 1'b0 ;
        reg_write_605 = 1'b0 ;
        reg_write_606 = 1'b0 ;
        reg_write_607 = 1'b0 ;
        reg_write_608 = 1'b0 ;
        reg_write_609 = 1'b0 ;
        reg_write_610 = 1'b0 ;
        reg_write_611 = 1'b0 ;
        reg_write_612 = 1'b0 ;
        reg_write_613 = 1'b0 ;
        reg_write_614 = 1'b0 ;
        reg_write_615 = 1'b0 ;
        reg_write_616 = 1'b0 ;
        reg_write_617 = 1'b0 ;
        reg_write_618 = 1'b0 ;
        reg_write_619 = 1'b0 ;
        reg_write_620 = 1'b0 ;
        reg_write_621 = 1'b0 ;
        reg_write_622 = 1'b0 ;
        reg_write_623 = 1'b0 ;
        reg_write_624 = 1'b0 ;
        reg_write_625 = 1'b0 ;
        reg_write_626 = 1'b0 ;
        reg_write_627 = 1'b0 ;
        reg_write_628 = 1'b0 ;
        reg_write_629 = 1'b0 ;
        reg_write_630 = 1'b0 ;
        reg_write_631 = 1'b0 ;
        reg_write_632 = 1'b0 ;
        reg_write_633 = 1'b0 ;
        reg_write_634 = 1'b0 ;
        reg_write_635 = 1'b0 ;
        reg_write_636 = 1'b0 ;
        reg_write_637 = 1'b0 ;
        reg_write_638 = 1'b0 ;
        reg_write_639 = 1'b0 ;
        reg_write_640 = 1'b0 ;
        reg_write_641 = 1'b0 ;
        reg_write_642 = 1'b0 ;
        reg_write_643 = 1'b0 ;
        reg_write_644 = 1'b0 ;
        reg_write_645 = 1'b0 ;
        reg_write_646 = 1'b0 ;
        reg_write_647 = 1'b0 ;
        reg_write_648 = 1'b0 ;
        reg_write_649 = 1'b0 ;
        reg_write_650 = 1'b0 ;
        reg_write_651 = 1'b0 ;
        reg_write_652 = 1'b0 ;
        reg_write_653 = 1'b0 ;
        reg_write_654 = 1'b0 ;
        reg_write_655 = 1'b0 ;
        reg_write_656 = 1'b0 ;
        reg_write_657 = 1'b0 ;
        reg_write_658 = 1'b0 ;
        reg_write_659 = 1'b0 ;
        reg_write_660 = 1'b0 ;
        reg_write_661 = 1'b0 ;
        reg_write_662 = 1'b0 ;
        reg_write_663 = 1'b0 ;
        reg_write_664 = 1'b0 ;
        reg_write_665 = 1'b0 ;
        reg_write_666 = 1'b0 ;
        reg_write_667 = 1'b0 ;
        reg_write_668 = 1'b0 ;
        reg_write_669 = 1'b0 ;
        reg_write_670 = 1'b0 ;
        reg_write_671 = 1'b0 ;
        reg_write_672 = 1'b0 ;
        reg_write_673 = 1'b0 ;
        reg_write_674 = 1'b0 ;
        reg_write_675 = 1'b0 ;
        reg_write_676 = 1'b0 ;
        reg_write_677 = 1'b0 ;
        reg_write_678 = 1'b0 ;
        reg_write_679 = 1'b0 ;
        reg_write_680 = 1'b0 ;
        reg_write_681 = 1'b0 ;
        reg_write_682 = 1'b0 ;
        reg_write_683 = 1'b0 ;
        reg_write_684 = 1'b0 ;
        reg_write_685 = 1'b0 ;
        reg_write_686 = 1'b0 ;
        reg_write_687 = 1'b0 ;
        reg_write_688 = 1'b0 ;
        reg_write_689 = 1'b0 ;
        reg_write_690 = 1'b0 ;
        reg_write_691 = 1'b0 ;
        reg_write_692 = 1'b0 ;
        reg_write_693 = 1'b0 ;
        reg_write_694 = 1'b0 ;
        reg_write_695 = 1'b0 ;
        reg_write_696 = 1'b0 ;
        reg_write_697 = 1'b0 ;
        reg_write_698 = 1'b0 ;
        reg_write_699 = 1'b0 ;
        reg_write_700 = 1'b0 ;
        reg_write_701 = 1'b0 ;
        reg_write_702 = 1'b0 ;
        reg_write_703 = 1'b0 ;
        reg_write_704 = 1'b0 ;
        reg_write_705 = 1'b0 ;
        reg_write_706 = 1'b0 ;
        reg_write_707 = 1'b0 ;
        reg_write_708 = 1'b0 ;
        reg_write_709 = 1'b0 ;
        reg_write_710 = 1'b0 ;
        reg_write_711 = 1'b0 ;
        reg_write_712 = 1'b0 ;
        reg_write_713 = 1'b0 ;
        reg_write_714 = 1'b0 ;
        reg_write_715 = 1'b0 ;
        reg_write_716 = 1'b0 ;
        reg_write_717 = 1'b0 ;
        reg_write_718 = 1'b0 ;
        reg_write_719 = 1'b0 ;
        reg_write_720 = 1'b0 ;
        reg_write_721 = 1'b0 ;
        reg_write_722 = 1'b0 ;
        reg_write_723 = 1'b0 ;
        reg_write_724 = 1'b0 ;
        reg_write_725 = 1'b0 ;
        reg_write_726 = 1'b0 ;
        reg_write_727 = 1'b0 ;
        reg_write_728 = 1'b0 ;
        reg_write_729 = 1'b0 ;
        reg_write_730 = 1'b0 ;
        reg_write_731 = 1'b0 ;
        reg_write_732 = 1'b0 ;
        reg_write_733 = 1'b0 ;
        reg_write_734 = 1'b0 ;
        reg_write_735 = 1'b0 ;
        reg_write_736 = 1'b0 ;
        reg_write_737 = 1'b0 ;
        reg_write_738 = 1'b0 ;
        reg_write_739 = 1'b0 ;
        reg_write_740 = 1'b0 ;
        reg_write_741 = 1'b0 ;
        reg_write_742 = 1'b0 ;
        reg_write_743 = 1'b0 ;
        reg_write_744 = 1'b0 ;
        reg_write_745 = 1'b0 ;
        reg_write_746 = 1'b0 ;
        reg_write_747 = 1'b0 ;
        reg_write_748 = 1'b0 ;
        reg_write_749 = 1'b0 ;
        reg_write_750 = 1'b0 ;
        reg_write_751 = 1'b0 ;
        reg_write_752 = 1'b0 ;
        reg_write_753 = 1'b0 ;
        reg_write_754 = 1'b0 ;
        reg_write_755 = 1'b0 ;
        reg_write_756 = 1'b0 ;
        reg_write_757 = 1'b0 ;
        reg_write_758 = 1'b0 ;
        reg_write_759 = 1'b0 ;
        reg_write_760 = 1'b0 ;
        reg_write_761 = 1'b0 ;
        reg_write_762 = 1'b0 ;
        reg_write_763 = 1'b0 ;
        reg_write_764 = 1'b0 ;
        reg_write_765 = 1'b0 ;
        reg_write_766 = 1'b0 ;
        reg_write_767 = 1'b0 ;
        reg_write_768 = 1'b0 ;
        reg_write_769 = 1'b0 ;
        reg_write_770 = 1'b0 ;
        reg_write_771 = 1'b0 ;
        reg_write_772 = 1'b0 ;
        reg_write_773 = 1'b0 ;
        reg_write_774 = 1'b0 ;
        reg_write_775 = 1'b0 ;
        reg_write_776 = 1'b0 ;
        reg_write_777 = 1'b0 ;
        reg_write_778 = 1'b0 ;
        reg_write_779 = 1'b0 ;
        reg_write_780 = 1'b0 ;
        reg_write_781 = 1'b0 ;
        reg_write_782 = 1'b0 ;
        reg_write_783 = 1'b0 ;
        reg_write_784 = 1'b0 ;
        reg_write_785 = 1'b0 ;
        reg_write_786 = 1'b0 ;
        reg_write_787 = 1'b0 ;
        reg_write_788 = 1'b0 ;
        reg_write_789 = 1'b0 ;
        reg_write_790 = 1'b0 ;
        reg_write_791 = 1'b0 ;
        reg_write_792 = 1'b0 ;
        reg_write_793 = 1'b0 ;
        reg_write_794 = 1'b0 ;
        reg_write_795 = 1'b0 ;
        reg_write_796 = 1'b0 ;
        reg_write_797 = 1'b0 ;
        reg_write_798 = 1'b0 ;
        reg_write_799 = 1'b0 ;
        reg_write_800 = 1'b0 ;
        reg_write_801 = 1'b0 ;
        reg_write_802 = 1'b0 ;
        reg_write_803 = 1'b0 ;
        reg_write_804 = 1'b0 ;
        reg_write_805 = 1'b0 ;
        reg_write_806 = 1'b0 ;
        reg_write_807 = 1'b0 ;
        reg_write_808 = 1'b0 ;
        reg_write_809 = 1'b0 ;
        reg_write_810 = 1'b0 ;
        reg_write_811 = 1'b0 ;
        reg_write_812 = 1'b0 ;
        reg_write_813 = 1'b0 ;
        reg_write_814 = 1'b0 ;
        reg_write_815 = 1'b0 ;
        reg_write_816 = 1'b0 ;
        reg_write_817 = 1'b0 ;
        reg_write_818 = 1'b0 ;
        reg_write_819 = 1'b0 ;
        reg_write_820 = 1'b0 ;
        reg_write_821 = 1'b0 ;
        reg_write_822 = 1'b0 ;
        reg_write_823 = 1'b0 ;
        reg_write_824 = 1'b0 ;
        reg_write_825 = 1'b0 ;
        reg_write_826 = 1'b0 ;
        reg_write_827 = 1'b0 ;
        reg_write_828 = 1'b0 ;
        reg_write_829 = 1'b0 ;
        reg_write_830 = 1'b0 ;
        reg_write_831 = 1'b0 ;
        reg_write_832 = 1'b0 ;
        reg_write_833 = 1'b0 ;
        reg_write_834 = 1'b0 ;
        reg_write_835 = 1'b0 ;
        reg_write_836 = 1'b0 ;
        reg_write_837 = 1'b0 ;
        reg_write_838 = 1'b0 ;
        reg_write_839 = 1'b0 ;
        reg_write_840 = 1'b0 ;
        reg_write_841 = 1'b0 ;
        reg_write_842 = 1'b0 ;
        reg_write_843 = 1'b0 ;
        reg_write_844 = 1'b0 ;
        reg_write_845 = 1'b0 ;
        reg_write_846 = 1'b0 ;
        reg_write_847 = 1'b0 ;
        reg_write_848 = 1'b0 ;
        reg_write_849 = 1'b0 ;
        reg_write_850 = 1'b0 ;
        reg_write_851 = 1'b0 ;
        reg_write_852 = 1'b0 ;
        reg_write_853 = 1'b0 ;
        reg_write_854 = 1'b0 ;
        reg_write_855 = 1'b0 ;
        reg_write_856 = 1'b0 ;
        reg_write_857 = 1'b0 ;
        reg_write_858 = 1'b0 ;
        reg_write_859 = 1'b0 ;
        reg_write_860 = 1'b0 ;
        reg_write_861 = 1'b0 ;
        reg_write_862 = 1'b0 ;
        reg_write_863 = 1'b0 ;
        reg_write_864 = 1'b0 ;
        reg_write_865 = 1'b0 ;
        reg_write_866 = 1'b0 ;
        reg_write_867 = 1'b0 ;
        reg_write_868 = 1'b0 ;
        reg_write_869 = 1'b0 ;
        reg_write_870 = 1'b0 ;
        reg_write_871 = 1'b0 ;
        reg_write_872 = 1'b0 ;
        reg_write_873 = 1'b0 ;
        reg_write_874 = 1'b0 ;
        reg_write_875 = 1'b0 ;
        reg_write_876 = 1'b0 ;
        reg_write_877 = 1'b0 ;
        reg_write_878 = 1'b0 ;
        reg_write_879 = 1'b0 ;
        reg_write_880 = 1'b0 ;
        reg_write_881 = 1'b0 ;
        reg_write_882 = 1'b0 ;
        reg_write_883 = 1'b0 ;
        reg_write_884 = 1'b0 ;
        reg_write_885 = 1'b0 ;
        reg_write_886 = 1'b0 ;
        reg_write_887 = 1'b0 ;
        reg_write_888 = 1'b0 ;
        reg_write_889 = 1'b0 ;
        reg_write_890 = 1'b0 ;
        reg_write_891 = 1'b0 ;
        reg_write_892 = 1'b0 ;
        reg_write_893 = 1'b0 ;
        reg_write_894 = 1'b0 ;
        reg_write_895 = 1'b0 ;
        reg_write_896 = 1'b0 ;
        reg_write_897 = 1'b0 ;
        reg_write_898 = 1'b0 ;
        reg_write_899 = 1'b0 ;
        reg_write_900 = 1'b0 ;
        reg_write_901 = 1'b0 ;
        reg_write_902 = 1'b0 ;
        reg_write_903 = 1'b0 ;
        reg_write_904 = 1'b0 ;
        reg_write_905 = 1'b0 ;
        reg_write_906 = 1'b0 ;
        reg_write_907 = 1'b0 ;
        reg_write_908 = 1'b0 ;
        reg_write_909 = 1'b0 ;
        reg_write_910 = 1'b0 ;
        reg_write_911 = 1'b0 ;
        reg_write_912 = 1'b0 ;
        reg_write_913 = 1'b0 ;
        reg_write_914 = 1'b0 ;
        reg_write_915 = 1'b0 ;
        reg_write_916 = 1'b0 ;
        reg_write_917 = 1'b0 ;
        reg_write_918 = 1'b0 ;
        reg_write_919 = 1'b0 ;
        reg_write_920 = 1'b0 ;
        reg_write_921 = 1'b0 ;
        reg_write_922 = 1'b0 ;
        reg_write_923 = 1'b0 ;
        reg_write_924 = 1'b0 ;
        reg_write_925 = 1'b0 ;
        reg_write_926 = 1'b0 ;
        reg_write_927 = 1'b0 ;
        reg_write_928 = 1'b0 ;
        reg_write_929 = 1'b0 ;
        reg_write_930 = 1'b0 ;
        reg_write_931 = 1'b0 ;
        reg_write_932 = 1'b0 ;
        reg_write_933 = 1'b0 ;
        reg_write_934 = 1'b0 ;
        reg_write_935 = 1'b0 ;
        reg_write_936 = 1'b0 ;
        reg_write_937 = 1'b0 ;
        reg_write_938 = 1'b0 ;
        reg_write_939 = 1'b0 ;
        reg_write_940 = 1'b0 ;
        reg_write_941 = 1'b0 ;
        reg_write_942 = 1'b0 ;
        reg_write_943 = 1'b0 ;
        reg_write_944 = 1'b0 ;
        reg_write_945 = 1'b0 ;
        reg_write_946 = 1'b0 ;
        reg_write_947 = 1'b0 ;
        reg_write_948 = 1'b0 ;
        reg_write_949 = 1'b0 ;
        reg_write_950 = 1'b0 ;
        reg_write_951 = 1'b0 ;
        reg_write_952 = 1'b0 ;
        reg_write_953 = 1'b0 ;
        reg_write_954 = 1'b0 ;
        reg_write_955 = 1'b0 ;
        reg_write_956 = 1'b0 ;
        reg_write_957 = 1'b0 ;
        reg_write_958 = 1'b0 ;
        reg_write_959 = 1'b0 ;
        reg_write_960 = 1'b0 ;
        reg_write_961 = 1'b0 ;
        reg_write_962 = 1'b0 ;
        reg_write_963 = 1'b0 ;
        reg_write_964 = 1'b0 ;
        reg_write_965 = 1'b0 ;
        reg_write_966 = 1'b0 ;
        reg_write_967 = 1'b0 ;
        reg_write_968 = 1'b0 ;
        reg_write_969 = 1'b0 ;
        reg_write_970 = 1'b0 ;
        reg_write_971 = 1'b0 ;
        reg_write_972 = 1'b0 ;
        reg_write_973 = 1'b0 ;
        reg_write_974 = 1'b0 ;
        reg_write_975 = 1'b0 ;
        reg_write_976 = 1'b0 ;
        reg_write_977 = 1'b0 ;
        reg_write_978 = 1'b0 ;
        reg_write_979 = 1'b0 ;
        reg_write_980 = 1'b0 ;
        reg_write_981 = 1'b0 ;
        reg_write_982 = 1'b0 ;
        reg_write_983 = 1'b0 ;
        reg_write_984 = 1'b0 ;
        reg_write_985 = 1'b0 ;
        reg_write_986 = 1'b0 ;
        reg_write_987 = 1'b0 ;
        reg_write_988 = 1'b0 ;
        reg_write_989 = 1'b0 ;
        reg_write_990 = 1'b0 ;
        reg_write_991 = 1'b0 ;
        reg_write_992 = 1'b0 ;
        reg_write_993 = 1'b0 ;
        reg_write_994 = 1'b0 ;
        reg_write_995 = 1'b0 ;
        reg_write_996 = 1'b0 ;
        reg_write_997 = 1'b0 ;
        reg_write_998 = 1'b0 ;
        reg_write_999 = 1'b0 ;
        reg_write_1000 = 1'b0 ;
			end
		end

endmodule
