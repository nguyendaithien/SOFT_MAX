`timescale 1 ns/10 ps
module LUT #(parameter DATA_WIDTH = 16 , DATA_WIDTH_OUT = 24) (
		data_in
	 ,data_out
);
	input [DATA_WIDTH-1:0] data_in;
	output reg [DATA_WIDTH_OUT-1:0] data_out;
always @(data_in) begin
	case(data_in) 	
    16'b1110110000000000 : data_out = 24'b000000000000000000110111;
    16'b1110110000000001 : data_out = 24'b000000000000000000110111;
    16'b1110110000000010 : data_out = 24'b000000000000000000110111;
    16'b1110110000000011 : data_out = 24'b000000000000000000110111;
    16'b1110110000000100 : data_out = 24'b000000000000000000110111;
    16'b1110110000000101 : data_out = 24'b000000000000000000110111;
    16'b1110110000000110 : data_out = 24'b000000000000000000110111;
    16'b1110110000000111 : data_out = 24'b000000000000000000110111;
    16'b1110110000001000 : data_out = 24'b000000000000000000110111;
    16'b1110110000001001 : data_out = 24'b000000000000000000110111;
    16'b1110110000001010 : data_out = 24'b000000000000000000110111;
    16'b1110110000001011 : data_out = 24'b000000000000000000110111;
    16'b1110110000001100 : data_out = 24'b000000000000000000110111;
    16'b1110110000001101 : data_out = 24'b000000000000000000110111;
    16'b1110110000001110 : data_out = 24'b000000000000000000110111;
    16'b1110110000001111 : data_out = 24'b000000000000000000111000;
    16'b1110110000010000 : data_out = 24'b000000000000000000111000;
    16'b1110110000010001 : data_out = 24'b000000000000000000111000;
    16'b1110110000010010 : data_out = 24'b000000000000000000111000;
    16'b1110110000010011 : data_out = 24'b000000000000000000111000;
    16'b1110110000010100 : data_out = 24'b000000000000000000111000;
    16'b1110110000010101 : data_out = 24'b000000000000000000111000;
    16'b1110110000010110 : data_out = 24'b000000000000000000111000;
    16'b1110110000010111 : data_out = 24'b000000000000000000111000;
    16'b1110110000011000 : data_out = 24'b000000000000000000111000;
    16'b1110110000011001 : data_out = 24'b000000000000000000111000;
    16'b1110110000011010 : data_out = 24'b000000000000000000111000;
    16'b1110110000011011 : data_out = 24'b000000000000000000111000;
    16'b1110110000011100 : data_out = 24'b000000000000000000111000;
    16'b1110110000011101 : data_out = 24'b000000000000000000111000;
    16'b1110110000011110 : data_out = 24'b000000000000000000111000;
    16'b1110110000011111 : data_out = 24'b000000000000000000111000;
    16'b1110110000100000 : data_out = 24'b000000000000000000111000;
    16'b1110110000100001 : data_out = 24'b000000000000000000111001;
    16'b1110110000100010 : data_out = 24'b000000000000000000111001;
    16'b1110110000100011 : data_out = 24'b000000000000000000111001;
    16'b1110110000100100 : data_out = 24'b000000000000000000111001;
    16'b1110110000100101 : data_out = 24'b000000000000000000111001;
    16'b1110110000100110 : data_out = 24'b000000000000000000111001;
    16'b1110110000100111 : data_out = 24'b000000000000000000111001;
    16'b1110110000101000 : data_out = 24'b000000000000000000111001;
    16'b1110110000101001 : data_out = 24'b000000000000000000111001;
    16'b1110110000101010 : data_out = 24'b000000000000000000111001;
    16'b1110110000101011 : data_out = 24'b000000000000000000111001;
    16'b1110110000101100 : data_out = 24'b000000000000000000111001;
    16'b1110110000101101 : data_out = 24'b000000000000000000111001;
    16'b1110110000101110 : data_out = 24'b000000000000000000111001;
    16'b1110110000101111 : data_out = 24'b000000000000000000111001;
    16'b1110110000110000 : data_out = 24'b000000000000000000111001;
    16'b1110110000110001 : data_out = 24'b000000000000000000111001;
    16'b1110110000110010 : data_out = 24'b000000000000000000111001;
    16'b1110110000110011 : data_out = 24'b000000000000000000111010;
    16'b1110110000110100 : data_out = 24'b000000000000000000111010;
    16'b1110110000110101 : data_out = 24'b000000000000000000111010;
    16'b1110110000110110 : data_out = 24'b000000000000000000111010;
    16'b1110110000110111 : data_out = 24'b000000000000000000111010;
    16'b1110110000111000 : data_out = 24'b000000000000000000111010;
    16'b1110110000111001 : data_out = 24'b000000000000000000111010;
    16'b1110110000111010 : data_out = 24'b000000000000000000111010;
    16'b1110110000111011 : data_out = 24'b000000000000000000111010;
    16'b1110110000111100 : data_out = 24'b000000000000000000111010;
    16'b1110110000111101 : data_out = 24'b000000000000000000111010;
    16'b1110110000111110 : data_out = 24'b000000000000000000111010;
    16'b1110110000111111 : data_out = 24'b000000000000000000111010;
    16'b1110110001000000 : data_out = 24'b000000000000000000111010;
    16'b1110110001000001 : data_out = 24'b000000000000000000111010;
    16'b1110110001000010 : data_out = 24'b000000000000000000111010;
    16'b1110110001000011 : data_out = 24'b000000000000000000111010;
    16'b1110110001000100 : data_out = 24'b000000000000000000111010;
    16'b1110110001000101 : data_out = 24'b000000000000000000111011;
    16'b1110110001000110 : data_out = 24'b000000000000000000111011;
    16'b1110110001000111 : data_out = 24'b000000000000000000111011;
    16'b1110110001001000 : data_out = 24'b000000000000000000111011;
    16'b1110110001001001 : data_out = 24'b000000000000000000111011;
    16'b1110110001001010 : data_out = 24'b000000000000000000111011;
    16'b1110110001001011 : data_out = 24'b000000000000000000111011;
    16'b1110110001001100 : data_out = 24'b000000000000000000111011;
    16'b1110110001001101 : data_out = 24'b000000000000000000111011;
    16'b1110110001001110 : data_out = 24'b000000000000000000111011;
    16'b1110110001001111 : data_out = 24'b000000000000000000111011;
    16'b1110110001010000 : data_out = 24'b000000000000000000111011;
    16'b1110110001010001 : data_out = 24'b000000000000000000111011;
    16'b1110110001010010 : data_out = 24'b000000000000000000111011;
    16'b1110110001010011 : data_out = 24'b000000000000000000111011;
    16'b1110110001010100 : data_out = 24'b000000000000000000111011;
    16'b1110110001010101 : data_out = 24'b000000000000000000111011;
    16'b1110110001010110 : data_out = 24'b000000000000000000111100;
    16'b1110110001010111 : data_out = 24'b000000000000000000111100;
    16'b1110110001011000 : data_out = 24'b000000000000000000111100;
    16'b1110110001011001 : data_out = 24'b000000000000000000111100;
    16'b1110110001011010 : data_out = 24'b000000000000000000111100;
    16'b1110110001011011 : data_out = 24'b000000000000000000111100;
    16'b1110110001011100 : data_out = 24'b000000000000000000111100;
    16'b1110110001011101 : data_out = 24'b000000000000000000111100;
    16'b1110110001011110 : data_out = 24'b000000000000000000111100;
    16'b1110110001011111 : data_out = 24'b000000000000000000111100;
    16'b1110110001100000 : data_out = 24'b000000000000000000111100;
    16'b1110110001100001 : data_out = 24'b000000000000000000111100;
    16'b1110110001100010 : data_out = 24'b000000000000000000111100;
    16'b1110110001100011 : data_out = 24'b000000000000000000111100;
    16'b1110110001100100 : data_out = 24'b000000000000000000111100;
    16'b1110110001100101 : data_out = 24'b000000000000000000111100;
    16'b1110110001100110 : data_out = 24'b000000000000000000111100;
    16'b1110110001100111 : data_out = 24'b000000000000000000111101;
    16'b1110110001101000 : data_out = 24'b000000000000000000111101;
    16'b1110110001101001 : data_out = 24'b000000000000000000111101;
    16'b1110110001101010 : data_out = 24'b000000000000000000111101;
    16'b1110110001101011 : data_out = 24'b000000000000000000111101;
    16'b1110110001101100 : data_out = 24'b000000000000000000111101;
    16'b1110110001101101 : data_out = 24'b000000000000000000111101;
    16'b1110110001101110 : data_out = 24'b000000000000000000111101;
    16'b1110110001101111 : data_out = 24'b000000000000000000111101;
    16'b1110110001110000 : data_out = 24'b000000000000000000111101;
    16'b1110110001110001 : data_out = 24'b000000000000000000111101;
    16'b1110110001110010 : data_out = 24'b000000000000000000111101;
    16'b1110110001110011 : data_out = 24'b000000000000000000111101;
    16'b1110110001110100 : data_out = 24'b000000000000000000111101;
    16'b1110110001110101 : data_out = 24'b000000000000000000111101;
    16'b1110110001110110 : data_out = 24'b000000000000000000111101;
    16'b1110110001110111 : data_out = 24'b000000000000000000111101;
    16'b1110110001111000 : data_out = 24'b000000000000000000111110;
    16'b1110110001111001 : data_out = 24'b000000000000000000111110;
    16'b1110110001111010 : data_out = 24'b000000000000000000111110;
    16'b1110110001111011 : data_out = 24'b000000000000000000111110;
    16'b1110110001111100 : data_out = 24'b000000000000000000111110;
    16'b1110110001111101 : data_out = 24'b000000000000000000111110;
    16'b1110110001111110 : data_out = 24'b000000000000000000111110;
    16'b1110110001111111 : data_out = 24'b000000000000000000111110;
    16'b1110110010000000 : data_out = 24'b000000000000000000111110;
    16'b1110110010000001 : data_out = 24'b000000000000000000111110;
    16'b1110110010000010 : data_out = 24'b000000000000000000111110;
    16'b1110110010000011 : data_out = 24'b000000000000000000111110;
    16'b1110110010000100 : data_out = 24'b000000000000000000111110;
    16'b1110110010000101 : data_out = 24'b000000000000000000111110;
    16'b1110110010000110 : data_out = 24'b000000000000000000111110;
    16'b1110110010000111 : data_out = 24'b000000000000000000111110;
    16'b1110110010001000 : data_out = 24'b000000000000000000111111;
    16'b1110110010001001 : data_out = 24'b000000000000000000111111;
    16'b1110110010001010 : data_out = 24'b000000000000000000111111;
    16'b1110110010001011 : data_out = 24'b000000000000000000111111;
    16'b1110110010001100 : data_out = 24'b000000000000000000111111;
    16'b1110110010001101 : data_out = 24'b000000000000000000111111;
    16'b1110110010001110 : data_out = 24'b000000000000000000111111;
    16'b1110110010001111 : data_out = 24'b000000000000000000111111;
    16'b1110110010010000 : data_out = 24'b000000000000000000111111;
    16'b1110110010010001 : data_out = 24'b000000000000000000111111;
    16'b1110110010010010 : data_out = 24'b000000000000000000111111;
    16'b1110110010010011 : data_out = 24'b000000000000000000111111;
    16'b1110110010010100 : data_out = 24'b000000000000000000111111;
    16'b1110110010010101 : data_out = 24'b000000000000000000111111;
    16'b1110110010010110 : data_out = 24'b000000000000000000111111;
    16'b1110110010010111 : data_out = 24'b000000000000000000111111;
    16'b1110110010011000 : data_out = 24'b000000000000000001000000;
    16'b1110110010011001 : data_out = 24'b000000000000000001000000;
    16'b1110110010011010 : data_out = 24'b000000000000000001000000;
    16'b1110110010011011 : data_out = 24'b000000000000000001000000;
    16'b1110110010011100 : data_out = 24'b000000000000000001000000;
    16'b1110110010011101 : data_out = 24'b000000000000000001000000;
    16'b1110110010011110 : data_out = 24'b000000000000000001000000;
    16'b1110110010011111 : data_out = 24'b000000000000000001000000;
    16'b1110110010100000 : data_out = 24'b000000000000000001000000;
    16'b1110110010100001 : data_out = 24'b000000000000000001000000;
    16'b1110110010100010 : data_out = 24'b000000000000000001000000;
    16'b1110110010100011 : data_out = 24'b000000000000000001000000;
    16'b1110110010100100 : data_out = 24'b000000000000000001000000;
    16'b1110110010100101 : data_out = 24'b000000000000000001000000;
    16'b1110110010100110 : data_out = 24'b000000000000000001000000;
    16'b1110110010100111 : data_out = 24'b000000000000000001000000;
    16'b1110110010101000 : data_out = 24'b000000000000000001000001;
    16'b1110110010101001 : data_out = 24'b000000000000000001000001;
    16'b1110110010101010 : data_out = 24'b000000000000000001000001;
    16'b1110110010101011 : data_out = 24'b000000000000000001000001;
    16'b1110110010101100 : data_out = 24'b000000000000000001000001;
    16'b1110110010101101 : data_out = 24'b000000000000000001000001;
    16'b1110110010101110 : data_out = 24'b000000000000000001000001;
    16'b1110110010101111 : data_out = 24'b000000000000000001000001;
    16'b1110110010110000 : data_out = 24'b000000000000000001000001;
    16'b1110110010110001 : data_out = 24'b000000000000000001000001;
    16'b1110110010110010 : data_out = 24'b000000000000000001000001;
    16'b1110110010110011 : data_out = 24'b000000000000000001000001;
    16'b1110110010110100 : data_out = 24'b000000000000000001000001;
    16'b1110110010110101 : data_out = 24'b000000000000000001000001;
    16'b1110110010110110 : data_out = 24'b000000000000000001000001;
    16'b1110110010110111 : data_out = 24'b000000000000000001000001;
    16'b1110110010111000 : data_out = 24'b000000000000000001000010;
    16'b1110110010111001 : data_out = 24'b000000000000000001000010;
    16'b1110110010111010 : data_out = 24'b000000000000000001000010;
    16'b1110110010111011 : data_out = 24'b000000000000000001000010;
    16'b1110110010111100 : data_out = 24'b000000000000000001000010;
    16'b1110110010111101 : data_out = 24'b000000000000000001000010;
    16'b1110110010111110 : data_out = 24'b000000000000000001000010;
    16'b1110110010111111 : data_out = 24'b000000000000000001000010;
    16'b1110110011000000 : data_out = 24'b000000000000000001000010;
    16'b1110110011000001 : data_out = 24'b000000000000000001000010;
    16'b1110110011000010 : data_out = 24'b000000000000000001000010;
    16'b1110110011000011 : data_out = 24'b000000000000000001000010;
    16'b1110110011000100 : data_out = 24'b000000000000000001000010;
    16'b1110110011000101 : data_out = 24'b000000000000000001000010;
    16'b1110110011000110 : data_out = 24'b000000000000000001000010;
    16'b1110110011000111 : data_out = 24'b000000000000000001000011;
    16'b1110110011001000 : data_out = 24'b000000000000000001000011;
    16'b1110110011001001 : data_out = 24'b000000000000000001000011;
    16'b1110110011001010 : data_out = 24'b000000000000000001000011;
    16'b1110110011001011 : data_out = 24'b000000000000000001000011;
    16'b1110110011001100 : data_out = 24'b000000000000000001000011;
    16'b1110110011001101 : data_out = 24'b000000000000000001000011;
    16'b1110110011001110 : data_out = 24'b000000000000000001000011;
    16'b1110110011001111 : data_out = 24'b000000000000000001000011;
    16'b1110110011010000 : data_out = 24'b000000000000000001000011;
    16'b1110110011010001 : data_out = 24'b000000000000000001000011;
    16'b1110110011010010 : data_out = 24'b000000000000000001000011;
    16'b1110110011010011 : data_out = 24'b000000000000000001000011;
    16'b1110110011010100 : data_out = 24'b000000000000000001000011;
    16'b1110110011010101 : data_out = 24'b000000000000000001000011;
    16'b1110110011010110 : data_out = 24'b000000000000000001000100;
    16'b1110110011010111 : data_out = 24'b000000000000000001000100;
    16'b1110110011011000 : data_out = 24'b000000000000000001000100;
    16'b1110110011011001 : data_out = 24'b000000000000000001000100;
    16'b1110110011011010 : data_out = 24'b000000000000000001000100;
    16'b1110110011011011 : data_out = 24'b000000000000000001000100;
    16'b1110110011011100 : data_out = 24'b000000000000000001000100;
    16'b1110110011011101 : data_out = 24'b000000000000000001000100;
    16'b1110110011011110 : data_out = 24'b000000000000000001000100;
    16'b1110110011011111 : data_out = 24'b000000000000000001000100;
    16'b1110110011100000 : data_out = 24'b000000000000000001000100;
    16'b1110110011100001 : data_out = 24'b000000000000000001000100;
    16'b1110110011100010 : data_out = 24'b000000000000000001000100;
    16'b1110110011100011 : data_out = 24'b000000000000000001000100;
    16'b1110110011100100 : data_out = 24'b000000000000000001000100;
    16'b1110110011100101 : data_out = 24'b000000000000000001000101;
    16'b1110110011100110 : data_out = 24'b000000000000000001000101;
    16'b1110110011100111 : data_out = 24'b000000000000000001000101;
    16'b1110110011101000 : data_out = 24'b000000000000000001000101;
    16'b1110110011101001 : data_out = 24'b000000000000000001000101;
    16'b1110110011101010 : data_out = 24'b000000000000000001000101;
    16'b1110110011101011 : data_out = 24'b000000000000000001000101;
    16'b1110110011101100 : data_out = 24'b000000000000000001000101;
    16'b1110110011101101 : data_out = 24'b000000000000000001000101;
    16'b1110110011101110 : data_out = 24'b000000000000000001000101;
    16'b1110110011101111 : data_out = 24'b000000000000000001000101;
    16'b1110110011110000 : data_out = 24'b000000000000000001000101;
    16'b1110110011110001 : data_out = 24'b000000000000000001000101;
    16'b1110110011110010 : data_out = 24'b000000000000000001000101;
    16'b1110110011110011 : data_out = 24'b000000000000000001000101;
    16'b1110110011110100 : data_out = 24'b000000000000000001000110;
    16'b1110110011110101 : data_out = 24'b000000000000000001000110;
    16'b1110110011110110 : data_out = 24'b000000000000000001000110;
    16'b1110110011110111 : data_out = 24'b000000000000000001000110;
    16'b1110110011111000 : data_out = 24'b000000000000000001000110;
    16'b1110110011111001 : data_out = 24'b000000000000000001000110;
    16'b1110110011111010 : data_out = 24'b000000000000000001000110;
    16'b1110110011111011 : data_out = 24'b000000000000000001000110;
    16'b1110110011111100 : data_out = 24'b000000000000000001000110;
    16'b1110110011111101 : data_out = 24'b000000000000000001000110;
    16'b1110110011111110 : data_out = 24'b000000000000000001000110;
    16'b1110110011111111 : data_out = 24'b000000000000000001000110;
    16'b1110110100000000 : data_out = 24'b000000000000000001000110;
    16'b1110110100000001 : data_out = 24'b000000000000000001000110;
    16'b1110110100000010 : data_out = 24'b000000000000000001000111;
    16'b1110110100000011 : data_out = 24'b000000000000000001000111;
    16'b1110110100000100 : data_out = 24'b000000000000000001000111;
    16'b1110110100000101 : data_out = 24'b000000000000000001000111;
    16'b1110110100000110 : data_out = 24'b000000000000000001000111;
    16'b1110110100000111 : data_out = 24'b000000000000000001000111;
    16'b1110110100001000 : data_out = 24'b000000000000000001000111;
    16'b1110110100001001 : data_out = 24'b000000000000000001000111;
    16'b1110110100001010 : data_out = 24'b000000000000000001000111;
    16'b1110110100001011 : data_out = 24'b000000000000000001000111;
    16'b1110110100001100 : data_out = 24'b000000000000000001000111;
    16'b1110110100001101 : data_out = 24'b000000000000000001000111;
    16'b1110110100001110 : data_out = 24'b000000000000000001000111;
    16'b1110110100001111 : data_out = 24'b000000000000000001000111;
    16'b1110110100010000 : data_out = 24'b000000000000000001000111;
    16'b1110110100010001 : data_out = 24'b000000000000000001001000;
    16'b1110110100010010 : data_out = 24'b000000000000000001001000;
    16'b1110110100010011 : data_out = 24'b000000000000000001001000;
    16'b1110110100010100 : data_out = 24'b000000000000000001001000;
    16'b1110110100010101 : data_out = 24'b000000000000000001001000;
    16'b1110110100010110 : data_out = 24'b000000000000000001001000;
    16'b1110110100010111 : data_out = 24'b000000000000000001001000;
    16'b1110110100011000 : data_out = 24'b000000000000000001001000;
    16'b1110110100011001 : data_out = 24'b000000000000000001001000;
    16'b1110110100011010 : data_out = 24'b000000000000000001001000;
    16'b1110110100011011 : data_out = 24'b000000000000000001001000;
    16'b1110110100011100 : data_out = 24'b000000000000000001001000;
    16'b1110110100011101 : data_out = 24'b000000000000000001001000;
    16'b1110110100011110 : data_out = 24'b000000000000000001001000;
    16'b1110110100011111 : data_out = 24'b000000000000000001001001;
    16'b1110110100100000 : data_out = 24'b000000000000000001001001;
    16'b1110110100100001 : data_out = 24'b000000000000000001001001;
    16'b1110110100100010 : data_out = 24'b000000000000000001001001;
    16'b1110110100100011 : data_out = 24'b000000000000000001001001;
    16'b1110110100100100 : data_out = 24'b000000000000000001001001;
    16'b1110110100100101 : data_out = 24'b000000000000000001001001;
    16'b1110110100100110 : data_out = 24'b000000000000000001001001;
    16'b1110110100100111 : data_out = 24'b000000000000000001001001;
    16'b1110110100101000 : data_out = 24'b000000000000000001001001;
    16'b1110110100101001 : data_out = 24'b000000000000000001001001;
    16'b1110110100101010 : data_out = 24'b000000000000000001001001;
    16'b1110110100101011 : data_out = 24'b000000000000000001001001;
    16'b1110110100101100 : data_out = 24'b000000000000000001001001;
    16'b1110110100101101 : data_out = 24'b000000000000000001001010;
    16'b1110110100101110 : data_out = 24'b000000000000000001001010;
    16'b1110110100101111 : data_out = 24'b000000000000000001001010;
    16'b1110110100110000 : data_out = 24'b000000000000000001001010;
    16'b1110110100110001 : data_out = 24'b000000000000000001001010;
    16'b1110110100110010 : data_out = 24'b000000000000000001001010;
    16'b1110110100110011 : data_out = 24'b000000000000000001001010;
    16'b1110110100110100 : data_out = 24'b000000000000000001001010;
    16'b1110110100110101 : data_out = 24'b000000000000000001001010;
    16'b1110110100110110 : data_out = 24'b000000000000000001001010;
    16'b1110110100110111 : data_out = 24'b000000000000000001001010;
    16'b1110110100111000 : data_out = 24'b000000000000000001001010;
    16'b1110110100111001 : data_out = 24'b000000000000000001001010;
    16'b1110110100111010 : data_out = 24'b000000000000000001001011;
    16'b1110110100111011 : data_out = 24'b000000000000000001001011;
    16'b1110110100111100 : data_out = 24'b000000000000000001001011;
    16'b1110110100111101 : data_out = 24'b000000000000000001001011;
    16'b1110110100111110 : data_out = 24'b000000000000000001001011;
    16'b1110110100111111 : data_out = 24'b000000000000000001001011;
    16'b1110110101000000 : data_out = 24'b000000000000000001001011;
    16'b1110110101000001 : data_out = 24'b000000000000000001001011;
    16'b1110110101000010 : data_out = 24'b000000000000000001001011;
    16'b1110110101000011 : data_out = 24'b000000000000000001001011;
    16'b1110110101000100 : data_out = 24'b000000000000000001001011;
    16'b1110110101000101 : data_out = 24'b000000000000000001001011;
    16'b1110110101000110 : data_out = 24'b000000000000000001001011;
    16'b1110110101000111 : data_out = 24'b000000000000000001001011;
    16'b1110110101001000 : data_out = 24'b000000000000000001001100;
    16'b1110110101001001 : data_out = 24'b000000000000000001001100;
    16'b1110110101001010 : data_out = 24'b000000000000000001001100;
    16'b1110110101001011 : data_out = 24'b000000000000000001001100;
    16'b1110110101001100 : data_out = 24'b000000000000000001001100;
    16'b1110110101001101 : data_out = 24'b000000000000000001001100;
    16'b1110110101001110 : data_out = 24'b000000000000000001001100;
    16'b1110110101001111 : data_out = 24'b000000000000000001001100;
    16'b1110110101010000 : data_out = 24'b000000000000000001001100;
    16'b1110110101010001 : data_out = 24'b000000000000000001001100;
    16'b1110110101010010 : data_out = 24'b000000000000000001001100;
    16'b1110110101010011 : data_out = 24'b000000000000000001001100;
    16'b1110110101010100 : data_out = 24'b000000000000000001001100;
    16'b1110110101010101 : data_out = 24'b000000000000000001001101;
    16'b1110110101010110 : data_out = 24'b000000000000000001001101;
    16'b1110110101010111 : data_out = 24'b000000000000000001001101;
    16'b1110110101011000 : data_out = 24'b000000000000000001001101;
    16'b1110110101011001 : data_out = 24'b000000000000000001001101;
    16'b1110110101011010 : data_out = 24'b000000000000000001001101;
    16'b1110110101011011 : data_out = 24'b000000000000000001001101;
    16'b1110110101011100 : data_out = 24'b000000000000000001001101;
    16'b1110110101011101 : data_out = 24'b000000000000000001001101;
    16'b1110110101011110 : data_out = 24'b000000000000000001001101;
    16'b1110110101011111 : data_out = 24'b000000000000000001001101;
    16'b1110110101100000 : data_out = 24'b000000000000000001001101;
    16'b1110110101100001 : data_out = 24'b000000000000000001001101;
    16'b1110110101100010 : data_out = 24'b000000000000000001001101;
    16'b1110110101100011 : data_out = 24'b000000000000000001001110;
    16'b1110110101100100 : data_out = 24'b000000000000000001001110;
    16'b1110110101100101 : data_out = 24'b000000000000000001001110;
    16'b1110110101100110 : data_out = 24'b000000000000000001001110;
    16'b1110110101100111 : data_out = 24'b000000000000000001001110;
    16'b1110110101101000 : data_out = 24'b000000000000000001001110;
    16'b1110110101101001 : data_out = 24'b000000000000000001001110;
    16'b1110110101101010 : data_out = 24'b000000000000000001001110;
    16'b1110110101101011 : data_out = 24'b000000000000000001001110;
    16'b1110110101101100 : data_out = 24'b000000000000000001001110;
    16'b1110110101101101 : data_out = 24'b000000000000000001001110;
    16'b1110110101101110 : data_out = 24'b000000000000000001001110;
    16'b1110110101101111 : data_out = 24'b000000000000000001001110;
    16'b1110110101110000 : data_out = 24'b000000000000000001001111;
    16'b1110110101110001 : data_out = 24'b000000000000000001001111;
    16'b1110110101110010 : data_out = 24'b000000000000000001001111;
    16'b1110110101110011 : data_out = 24'b000000000000000001001111;
    16'b1110110101110100 : data_out = 24'b000000000000000001001111;
    16'b1110110101110101 : data_out = 24'b000000000000000001001111;
    16'b1110110101110110 : data_out = 24'b000000000000000001001111;
    16'b1110110101110111 : data_out = 24'b000000000000000001001111;
    16'b1110110101111000 : data_out = 24'b000000000000000001001111;
    16'b1110110101111001 : data_out = 24'b000000000000000001001111;
    16'b1110110101111010 : data_out = 24'b000000000000000001001111;
    16'b1110110101111011 : data_out = 24'b000000000000000001001111;
    16'b1110110101111100 : data_out = 24'b000000000000000001001111;
    16'b1110110101111101 : data_out = 24'b000000000000000001010000;
    16'b1110110101111110 : data_out = 24'b000000000000000001010000;
    16'b1110110101111111 : data_out = 24'b000000000000000001010000;
    16'b1110110110000000 : data_out = 24'b000000000000000001010000;
    16'b1110110110000001 : data_out = 24'b000000000000000001010000;
    16'b1110110110000010 : data_out = 24'b000000000000000001010000;
    16'b1110110110000011 : data_out = 24'b000000000000000001010000;
    16'b1110110110000100 : data_out = 24'b000000000000000001010000;
    16'b1110110110000101 : data_out = 24'b000000000000000001010000;
    16'b1110110110000110 : data_out = 24'b000000000000000001010000;
    16'b1110110110000111 : data_out = 24'b000000000000000001010000;
    16'b1110110110001000 : data_out = 24'b000000000000000001010000;
    16'b1110110110001001 : data_out = 24'b000000000000000001010001;
    16'b1110110110001010 : data_out = 24'b000000000000000001010001;
    16'b1110110110001011 : data_out = 24'b000000000000000001010001;
    16'b1110110110001100 : data_out = 24'b000000000000000001010001;
    16'b1110110110001101 : data_out = 24'b000000000000000001010001;
    16'b1110110110001110 : data_out = 24'b000000000000000001010001;
    16'b1110110110001111 : data_out = 24'b000000000000000001010001;
    16'b1110110110010000 : data_out = 24'b000000000000000001010001;
    16'b1110110110010001 : data_out = 24'b000000000000000001010001;
    16'b1110110110010010 : data_out = 24'b000000000000000001010001;
    16'b1110110110010011 : data_out = 24'b000000000000000001010001;
    16'b1110110110010100 : data_out = 24'b000000000000000001010001;
    16'b1110110110010101 : data_out = 24'b000000000000000001010001;
    16'b1110110110010110 : data_out = 24'b000000000000000001010010;
    16'b1110110110010111 : data_out = 24'b000000000000000001010010;
    16'b1110110110011000 : data_out = 24'b000000000000000001010010;
    16'b1110110110011001 : data_out = 24'b000000000000000001010010;
    16'b1110110110011010 : data_out = 24'b000000000000000001010010;
    16'b1110110110011011 : data_out = 24'b000000000000000001010010;
    16'b1110110110011100 : data_out = 24'b000000000000000001010010;
    16'b1110110110011101 : data_out = 24'b000000000000000001010010;
    16'b1110110110011110 : data_out = 24'b000000000000000001010010;
    16'b1110110110011111 : data_out = 24'b000000000000000001010010;
    16'b1110110110100000 : data_out = 24'b000000000000000001010010;
    16'b1110110110100001 : data_out = 24'b000000000000000001010010;
    16'b1110110110100010 : data_out = 24'b000000000000000001010011;
    16'b1110110110100011 : data_out = 24'b000000000000000001010011;
    16'b1110110110100100 : data_out = 24'b000000000000000001010011;
    16'b1110110110100101 : data_out = 24'b000000000000000001010011;
    16'b1110110110100110 : data_out = 24'b000000000000000001010011;
    16'b1110110110100111 : data_out = 24'b000000000000000001010011;
    16'b1110110110101000 : data_out = 24'b000000000000000001010011;
    16'b1110110110101001 : data_out = 24'b000000000000000001010011;
    16'b1110110110101010 : data_out = 24'b000000000000000001010011;
    16'b1110110110101011 : data_out = 24'b000000000000000001010011;
    16'b1110110110101100 : data_out = 24'b000000000000000001010011;
    16'b1110110110101101 : data_out = 24'b000000000000000001010011;
    16'b1110110110101110 : data_out = 24'b000000000000000001010100;
    16'b1110110110101111 : data_out = 24'b000000000000000001010100;
    16'b1110110110110000 : data_out = 24'b000000000000000001010100;
    16'b1110110110110001 : data_out = 24'b000000000000000001010100;
    16'b1110110110110010 : data_out = 24'b000000000000000001010100;
    16'b1110110110110011 : data_out = 24'b000000000000000001010100;
    16'b1110110110110100 : data_out = 24'b000000000000000001010100;
    16'b1110110110110101 : data_out = 24'b000000000000000001010100;
    16'b1110110110110110 : data_out = 24'b000000000000000001010100;
    16'b1110110110110111 : data_out = 24'b000000000000000001010100;
    16'b1110110110111000 : data_out = 24'b000000000000000001010100;
    16'b1110110110111001 : data_out = 24'b000000000000000001010100;
    16'b1110110110111010 : data_out = 24'b000000000000000001010100;
    16'b1110110110111011 : data_out = 24'b000000000000000001010101;
    16'b1110110110111100 : data_out = 24'b000000000000000001010101;
    16'b1110110110111101 : data_out = 24'b000000000000000001010101;
    16'b1110110110111110 : data_out = 24'b000000000000000001010101;
    16'b1110110110111111 : data_out = 24'b000000000000000001010101;
    16'b1110110111000000 : data_out = 24'b000000000000000001010101;
    16'b1110110111000001 : data_out = 24'b000000000000000001010101;
    16'b1110110111000010 : data_out = 24'b000000000000000001010101;
    16'b1110110111000011 : data_out = 24'b000000000000000001010101;
    16'b1110110111000100 : data_out = 24'b000000000000000001010101;
    16'b1110110111000101 : data_out = 24'b000000000000000001010101;
    16'b1110110111000110 : data_out = 24'b000000000000000001010101;
    16'b1110110111000111 : data_out = 24'b000000000000000001010110;
    16'b1110110111001000 : data_out = 24'b000000000000000001010110;
    16'b1110110111001001 : data_out = 24'b000000000000000001010110;
    16'b1110110111001010 : data_out = 24'b000000000000000001010110;
    16'b1110110111001011 : data_out = 24'b000000000000000001010110;
    16'b1110110111001100 : data_out = 24'b000000000000000001010110;
    16'b1110110111001101 : data_out = 24'b000000000000000001010110;
    16'b1110110111001110 : data_out = 24'b000000000000000001010110;
    16'b1110110111001111 : data_out = 24'b000000000000000001010110;
    16'b1110110111010000 : data_out = 24'b000000000000000001010110;
    16'b1110110111010001 : data_out = 24'b000000000000000001010110;
    16'b1110110111010010 : data_out = 24'b000000000000000001010111;
    16'b1110110111010011 : data_out = 24'b000000000000000001010111;
    16'b1110110111010100 : data_out = 24'b000000000000000001010111;
    16'b1110110111010101 : data_out = 24'b000000000000000001010111;
    16'b1110110111010110 : data_out = 24'b000000000000000001010111;
    16'b1110110111010111 : data_out = 24'b000000000000000001010111;
    16'b1110110111011000 : data_out = 24'b000000000000000001010111;
    16'b1110110111011001 : data_out = 24'b000000000000000001010111;
    16'b1110110111011010 : data_out = 24'b000000000000000001010111;
    16'b1110110111011011 : data_out = 24'b000000000000000001010111;
    16'b1110110111011100 : data_out = 24'b000000000000000001010111;
    16'b1110110111011101 : data_out = 24'b000000000000000001010111;
    16'b1110110111011110 : data_out = 24'b000000000000000001011000;
    16'b1110110111011111 : data_out = 24'b000000000000000001011000;
    16'b1110110111100000 : data_out = 24'b000000000000000001011000;
    16'b1110110111100001 : data_out = 24'b000000000000000001011000;
    16'b1110110111100010 : data_out = 24'b000000000000000001011000;
    16'b1110110111100011 : data_out = 24'b000000000000000001011000;
    16'b1110110111100100 : data_out = 24'b000000000000000001011000;
    16'b1110110111100101 : data_out = 24'b000000000000000001011000;
    16'b1110110111100110 : data_out = 24'b000000000000000001011000;
    16'b1110110111100111 : data_out = 24'b000000000000000001011000;
    16'b1110110111101000 : data_out = 24'b000000000000000001011000;
    16'b1110110111101001 : data_out = 24'b000000000000000001011000;
    16'b1110110111101010 : data_out = 24'b000000000000000001011001;
    16'b1110110111101011 : data_out = 24'b000000000000000001011001;
    16'b1110110111101100 : data_out = 24'b000000000000000001011001;
    16'b1110110111101101 : data_out = 24'b000000000000000001011001;
    16'b1110110111101110 : data_out = 24'b000000000000000001011001;
    16'b1110110111101111 : data_out = 24'b000000000000000001011001;
    16'b1110110111110000 : data_out = 24'b000000000000000001011001;
    16'b1110110111110001 : data_out = 24'b000000000000000001011001;
    16'b1110110111110010 : data_out = 24'b000000000000000001011001;
    16'b1110110111110011 : data_out = 24'b000000000000000001011001;
    16'b1110110111110100 : data_out = 24'b000000000000000001011001;
    16'b1110110111110101 : data_out = 24'b000000000000000001011010;
    16'b1110110111110110 : data_out = 24'b000000000000000001011010;
    16'b1110110111110111 : data_out = 24'b000000000000000001011010;
    16'b1110110111111000 : data_out = 24'b000000000000000001011010;
    16'b1110110111111001 : data_out = 24'b000000000000000001011010;
    16'b1110110111111010 : data_out = 24'b000000000000000001011010;
    16'b1110110111111011 : data_out = 24'b000000000000000001011010;
    16'b1110110111111100 : data_out = 24'b000000000000000001011010;
    16'b1110110111111101 : data_out = 24'b000000000000000001011010;
    16'b1110110111111110 : data_out = 24'b000000000000000001011010;
    16'b1110110111111111 : data_out = 24'b000000000000000001011010;
    16'b1110111000000000 : data_out = 24'b000000000000000001011011;
    16'b1110111000000001 : data_out = 24'b000000000000000001011011;
    16'b1110111000000010 : data_out = 24'b000000000000000001011011;
    16'b1110111000000011 : data_out = 24'b000000000000000001011011;
    16'b1110111000000100 : data_out = 24'b000000000000000001011011;
    16'b1110111000000101 : data_out = 24'b000000000000000001011011;
    16'b1110111000000110 : data_out = 24'b000000000000000001011011;
    16'b1110111000000111 : data_out = 24'b000000000000000001011011;
    16'b1110111000001000 : data_out = 24'b000000000000000001011011;
    16'b1110111000001001 : data_out = 24'b000000000000000001011011;
    16'b1110111000001010 : data_out = 24'b000000000000000001011011;
    16'b1110111000001011 : data_out = 24'b000000000000000001011011;
    16'b1110111000001100 : data_out = 24'b000000000000000001011100;
    16'b1110111000001101 : data_out = 24'b000000000000000001011100;
    16'b1110111000001110 : data_out = 24'b000000000000000001011100;
    16'b1110111000001111 : data_out = 24'b000000000000000001011100;
    16'b1110111000010000 : data_out = 24'b000000000000000001011100;
    16'b1110111000010001 : data_out = 24'b000000000000000001011100;
    16'b1110111000010010 : data_out = 24'b000000000000000001011100;
    16'b1110111000010011 : data_out = 24'b000000000000000001011100;
    16'b1110111000010100 : data_out = 24'b000000000000000001011100;
    16'b1110111000010101 : data_out = 24'b000000000000000001011100;
    16'b1110111000010110 : data_out = 24'b000000000000000001011100;
    16'b1110111000010111 : data_out = 24'b000000000000000001011101;
    16'b1110111000011000 : data_out = 24'b000000000000000001011101;
    16'b1110111000011001 : data_out = 24'b000000000000000001011101;
    16'b1110111000011010 : data_out = 24'b000000000000000001011101;
    16'b1110111000011011 : data_out = 24'b000000000000000001011101;
    16'b1110111000011100 : data_out = 24'b000000000000000001011101;
    16'b1110111000011101 : data_out = 24'b000000000000000001011101;
    16'b1110111000011110 : data_out = 24'b000000000000000001011101;
    16'b1110111000011111 : data_out = 24'b000000000000000001011101;
    16'b1110111000100000 : data_out = 24'b000000000000000001011101;
    16'b1110111000100001 : data_out = 24'b000000000000000001011101;
    16'b1110111000100010 : data_out = 24'b000000000000000001011110;
    16'b1110111000100011 : data_out = 24'b000000000000000001011110;
    16'b1110111000100100 : data_out = 24'b000000000000000001011110;
    16'b1110111000100101 : data_out = 24'b000000000000000001011110;
    16'b1110111000100110 : data_out = 24'b000000000000000001011110;
    16'b1110111000100111 : data_out = 24'b000000000000000001011110;
    16'b1110111000101000 : data_out = 24'b000000000000000001011110;
    16'b1110111000101001 : data_out = 24'b000000000000000001011110;
    16'b1110111000101010 : data_out = 24'b000000000000000001011110;
    16'b1110111000101011 : data_out = 24'b000000000000000001011110;
    16'b1110111000101100 : data_out = 24'b000000000000000001011111;
    16'b1110111000101101 : data_out = 24'b000000000000000001011111;
    16'b1110111000101110 : data_out = 24'b000000000000000001011111;
    16'b1110111000101111 : data_out = 24'b000000000000000001011111;
    16'b1110111000110000 : data_out = 24'b000000000000000001011111;
    16'b1110111000110001 : data_out = 24'b000000000000000001011111;
    16'b1110111000110010 : data_out = 24'b000000000000000001011111;
    16'b1110111000110011 : data_out = 24'b000000000000000001011111;
    16'b1110111000110100 : data_out = 24'b000000000000000001011111;
    16'b1110111000110101 : data_out = 24'b000000000000000001011111;
    16'b1110111000110110 : data_out = 24'b000000000000000001011111;
    16'b1110111000110111 : data_out = 24'b000000000000000001100000;
    16'b1110111000111000 : data_out = 24'b000000000000000001100000;
    16'b1110111000111001 : data_out = 24'b000000000000000001100000;
    16'b1110111000111010 : data_out = 24'b000000000000000001100000;
    16'b1110111000111011 : data_out = 24'b000000000000000001100000;
    16'b1110111000111100 : data_out = 24'b000000000000000001100000;
    16'b1110111000111101 : data_out = 24'b000000000000000001100000;
    16'b1110111000111110 : data_out = 24'b000000000000000001100000;
    16'b1110111000111111 : data_out = 24'b000000000000000001100000;
    16'b1110111001000000 : data_out = 24'b000000000000000001100000;
    16'b1110111001000001 : data_out = 24'b000000000000000001100000;
    16'b1110111001000010 : data_out = 24'b000000000000000001100001;
    16'b1110111001000011 : data_out = 24'b000000000000000001100001;
    16'b1110111001000100 : data_out = 24'b000000000000000001100001;
    16'b1110111001000101 : data_out = 24'b000000000000000001100001;
    16'b1110111001000110 : data_out = 24'b000000000000000001100001;
    16'b1110111001000111 : data_out = 24'b000000000000000001100001;
    16'b1110111001001000 : data_out = 24'b000000000000000001100001;
    16'b1110111001001001 : data_out = 24'b000000000000000001100001;
    16'b1110111001001010 : data_out = 24'b000000000000000001100001;
    16'b1110111001001011 : data_out = 24'b000000000000000001100001;
    16'b1110111001001100 : data_out = 24'b000000000000000001100010;
    16'b1110111001001101 : data_out = 24'b000000000000000001100010;
    16'b1110111001001110 : data_out = 24'b000000000000000001100010;
    16'b1110111001001111 : data_out = 24'b000000000000000001100010;
    16'b1110111001010000 : data_out = 24'b000000000000000001100010;
    16'b1110111001010001 : data_out = 24'b000000000000000001100010;
    16'b1110111001010010 : data_out = 24'b000000000000000001100010;
    16'b1110111001010011 : data_out = 24'b000000000000000001100010;
    16'b1110111001010100 : data_out = 24'b000000000000000001100010;
    16'b1110111001010101 : data_out = 24'b000000000000000001100010;
    16'b1110111001010110 : data_out = 24'b000000000000000001100010;
    16'b1110111001010111 : data_out = 24'b000000000000000001100011;
    16'b1110111001011000 : data_out = 24'b000000000000000001100011;
    16'b1110111001011001 : data_out = 24'b000000000000000001100011;
    16'b1110111001011010 : data_out = 24'b000000000000000001100011;
    16'b1110111001011011 : data_out = 24'b000000000000000001100011;
    16'b1110111001011100 : data_out = 24'b000000000000000001100011;
    16'b1110111001011101 : data_out = 24'b000000000000000001100011;
    16'b1110111001011110 : data_out = 24'b000000000000000001100011;
    16'b1110111001011111 : data_out = 24'b000000000000000001100011;
    16'b1110111001100000 : data_out = 24'b000000000000000001100011;
    16'b1110111001100001 : data_out = 24'b000000000000000001100100;
    16'b1110111001100010 : data_out = 24'b000000000000000001100100;
    16'b1110111001100011 : data_out = 24'b000000000000000001100100;
    16'b1110111001100100 : data_out = 24'b000000000000000001100100;
    16'b1110111001100101 : data_out = 24'b000000000000000001100100;
    16'b1110111001100110 : data_out = 24'b000000000000000001100100;
    16'b1110111001100111 : data_out = 24'b000000000000000001100100;
    16'b1110111001101000 : data_out = 24'b000000000000000001100100;
    16'b1110111001101001 : data_out = 24'b000000000000000001100100;
    16'b1110111001101010 : data_out = 24'b000000000000000001100100;
    16'b1110111001101011 : data_out = 24'b000000000000000001100101;
    16'b1110111001101100 : data_out = 24'b000000000000000001100101;
    16'b1110111001101101 : data_out = 24'b000000000000000001100101;
    16'b1110111001101110 : data_out = 24'b000000000000000001100101;
    16'b1110111001101111 : data_out = 24'b000000000000000001100101;
    16'b1110111001110000 : data_out = 24'b000000000000000001100101;
    16'b1110111001110001 : data_out = 24'b000000000000000001100101;
    16'b1110111001110010 : data_out = 24'b000000000000000001100101;
    16'b1110111001110011 : data_out = 24'b000000000000000001100101;
    16'b1110111001110100 : data_out = 24'b000000000000000001100101;
    16'b1110111001110101 : data_out = 24'b000000000000000001100110;
    16'b1110111001110110 : data_out = 24'b000000000000000001100110;
    16'b1110111001110111 : data_out = 24'b000000000000000001100110;
    16'b1110111001111000 : data_out = 24'b000000000000000001100110;
    16'b1110111001111001 : data_out = 24'b000000000000000001100110;
    16'b1110111001111010 : data_out = 24'b000000000000000001100110;
    16'b1110111001111011 : data_out = 24'b000000000000000001100110;
    16'b1110111001111100 : data_out = 24'b000000000000000001100110;
    16'b1110111001111101 : data_out = 24'b000000000000000001100110;
    16'b1110111001111110 : data_out = 24'b000000000000000001100110;
    16'b1110111001111111 : data_out = 24'b000000000000000001100111;
    16'b1110111010000000 : data_out = 24'b000000000000000001100111;
    16'b1110111010000001 : data_out = 24'b000000000000000001100111;
    16'b1110111010000010 : data_out = 24'b000000000000000001100111;
    16'b1110111010000011 : data_out = 24'b000000000000000001100111;
    16'b1110111010000100 : data_out = 24'b000000000000000001100111;
    16'b1110111010000101 : data_out = 24'b000000000000000001100111;
    16'b1110111010000110 : data_out = 24'b000000000000000001100111;
    16'b1110111010000111 : data_out = 24'b000000000000000001100111;
    16'b1110111010001000 : data_out = 24'b000000000000000001100111;
    16'b1110111010001001 : data_out = 24'b000000000000000001101000;
    16'b1110111010001010 : data_out = 24'b000000000000000001101000;
    16'b1110111010001011 : data_out = 24'b000000000000000001101000;
    16'b1110111010001100 : data_out = 24'b000000000000000001101000;
    16'b1110111010001101 : data_out = 24'b000000000000000001101000;
    16'b1110111010001110 : data_out = 24'b000000000000000001101000;
    16'b1110111010001111 : data_out = 24'b000000000000000001101000;
    16'b1110111010010000 : data_out = 24'b000000000000000001101000;
    16'b1110111010010001 : data_out = 24'b000000000000000001101000;
    16'b1110111010010010 : data_out = 24'b000000000000000001101000;
    16'b1110111010010011 : data_out = 24'b000000000000000001101001;
    16'b1110111010010100 : data_out = 24'b000000000000000001101001;
    16'b1110111010010101 : data_out = 24'b000000000000000001101001;
    16'b1110111010010110 : data_out = 24'b000000000000000001101001;
    16'b1110111010010111 : data_out = 24'b000000000000000001101001;
    16'b1110111010011000 : data_out = 24'b000000000000000001101001;
    16'b1110111010011001 : data_out = 24'b000000000000000001101001;
    16'b1110111010011010 : data_out = 24'b000000000000000001101001;
    16'b1110111010011011 : data_out = 24'b000000000000000001101001;
    16'b1110111010011100 : data_out = 24'b000000000000000001101001;
    16'b1110111010011101 : data_out = 24'b000000000000000001101010;
    16'b1110111010011110 : data_out = 24'b000000000000000001101010;
    16'b1110111010011111 : data_out = 24'b000000000000000001101010;
    16'b1110111010100000 : data_out = 24'b000000000000000001101010;
    16'b1110111010100001 : data_out = 24'b000000000000000001101010;
    16'b1110111010100010 : data_out = 24'b000000000000000001101010;
    16'b1110111010100011 : data_out = 24'b000000000000000001101010;
    16'b1110111010100100 : data_out = 24'b000000000000000001101010;
    16'b1110111010100101 : data_out = 24'b000000000000000001101010;
    16'b1110111010100110 : data_out = 24'b000000000000000001101011;
    16'b1110111010100111 : data_out = 24'b000000000000000001101011;
    16'b1110111010101000 : data_out = 24'b000000000000000001101011;
    16'b1110111010101001 : data_out = 24'b000000000000000001101011;
    16'b1110111010101010 : data_out = 24'b000000000000000001101011;
    16'b1110111010101011 : data_out = 24'b000000000000000001101011;
    16'b1110111010101100 : data_out = 24'b000000000000000001101011;
    16'b1110111010101101 : data_out = 24'b000000000000000001101011;
    16'b1110111010101110 : data_out = 24'b000000000000000001101011;
    16'b1110111010101111 : data_out = 24'b000000000000000001101011;
    16'b1110111010110000 : data_out = 24'b000000000000000001101100;
    16'b1110111010110001 : data_out = 24'b000000000000000001101100;
    16'b1110111010110010 : data_out = 24'b000000000000000001101100;
    16'b1110111010110011 : data_out = 24'b000000000000000001101100;
    16'b1110111010110100 : data_out = 24'b000000000000000001101100;
    16'b1110111010110101 : data_out = 24'b000000000000000001101100;
    16'b1110111010110110 : data_out = 24'b000000000000000001101100;
    16'b1110111010110111 : data_out = 24'b000000000000000001101100;
    16'b1110111010111000 : data_out = 24'b000000000000000001101100;
    16'b1110111010111001 : data_out = 24'b000000000000000001101101;
    16'b1110111010111010 : data_out = 24'b000000000000000001101101;
    16'b1110111010111011 : data_out = 24'b000000000000000001101101;
    16'b1110111010111100 : data_out = 24'b000000000000000001101101;
    16'b1110111010111101 : data_out = 24'b000000000000000001101101;
    16'b1110111010111110 : data_out = 24'b000000000000000001101101;
    16'b1110111010111111 : data_out = 24'b000000000000000001101101;
    16'b1110111011000000 : data_out = 24'b000000000000000001101101;
    16'b1110111011000001 : data_out = 24'b000000000000000001101101;
    16'b1110111011000010 : data_out = 24'b000000000000000001101101;
    16'b1110111011000011 : data_out = 24'b000000000000000001101110;
    16'b1110111011000100 : data_out = 24'b000000000000000001101110;
    16'b1110111011000101 : data_out = 24'b000000000000000001101110;
    16'b1110111011000110 : data_out = 24'b000000000000000001101110;
    16'b1110111011000111 : data_out = 24'b000000000000000001101110;
    16'b1110111011001000 : data_out = 24'b000000000000000001101110;
    16'b1110111011001001 : data_out = 24'b000000000000000001101110;
    16'b1110111011001010 : data_out = 24'b000000000000000001101110;
    16'b1110111011001011 : data_out = 24'b000000000000000001101110;
    16'b1110111011001100 : data_out = 24'b000000000000000001101111;
    16'b1110111011001101 : data_out = 24'b000000000000000001101111;
    16'b1110111011001110 : data_out = 24'b000000000000000001101111;
    16'b1110111011001111 : data_out = 24'b000000000000000001101111;
    16'b1110111011010000 : data_out = 24'b000000000000000001101111;
    16'b1110111011010001 : data_out = 24'b000000000000000001101111;
    16'b1110111011010010 : data_out = 24'b000000000000000001101111;
    16'b1110111011010011 : data_out = 24'b000000000000000001101111;
    16'b1110111011010100 : data_out = 24'b000000000000000001101111;
    16'b1110111011010101 : data_out = 24'b000000000000000001110000;
    16'b1110111011010110 : data_out = 24'b000000000000000001110000;
    16'b1110111011010111 : data_out = 24'b000000000000000001110000;
    16'b1110111011011000 : data_out = 24'b000000000000000001110000;
    16'b1110111011011001 : data_out = 24'b000000000000000001110000;
    16'b1110111011011010 : data_out = 24'b000000000000000001110000;
    16'b1110111011011011 : data_out = 24'b000000000000000001110000;
    16'b1110111011011100 : data_out = 24'b000000000000000001110000;
    16'b1110111011011101 : data_out = 24'b000000000000000001110000;
    16'b1110111011011110 : data_out = 24'b000000000000000001110001;
    16'b1110111011011111 : data_out = 24'b000000000000000001110001;
    16'b1110111011100000 : data_out = 24'b000000000000000001110001;
    16'b1110111011100001 : data_out = 24'b000000000000000001110001;
    16'b1110111011100010 : data_out = 24'b000000000000000001110001;
    16'b1110111011100011 : data_out = 24'b000000000000000001110001;
    16'b1110111011100100 : data_out = 24'b000000000000000001110001;
    16'b1110111011100101 : data_out = 24'b000000000000000001110001;
    16'b1110111011100110 : data_out = 24'b000000000000000001110001;
    16'b1110111011100111 : data_out = 24'b000000000000000001110010;
    16'b1110111011101000 : data_out = 24'b000000000000000001110010;
    16'b1110111011101001 : data_out = 24'b000000000000000001110010;
    16'b1110111011101010 : data_out = 24'b000000000000000001110010;
    16'b1110111011101011 : data_out = 24'b000000000000000001110010;
    16'b1110111011101100 : data_out = 24'b000000000000000001110010;
    16'b1110111011101101 : data_out = 24'b000000000000000001110010;
    16'b1110111011101110 : data_out = 24'b000000000000000001110010;
    16'b1110111011101111 : data_out = 24'b000000000000000001110010;
    16'b1110111011110000 : data_out = 24'b000000000000000001110011;
    16'b1110111011110001 : data_out = 24'b000000000000000001110011;
    16'b1110111011110010 : data_out = 24'b000000000000000001110011;
    16'b1110111011110011 : data_out = 24'b000000000000000001110011;
    16'b1110111011110100 : data_out = 24'b000000000000000001110011;
    16'b1110111011110101 : data_out = 24'b000000000000000001110011;
    16'b1110111011110110 : data_out = 24'b000000000000000001110011;
    16'b1110111011110111 : data_out = 24'b000000000000000001110011;
    16'b1110111011111000 : data_out = 24'b000000000000000001110011;
    16'b1110111011111001 : data_out = 24'b000000000000000001110100;
    16'b1110111011111010 : data_out = 24'b000000000000000001110100;
    16'b1110111011111011 : data_out = 24'b000000000000000001110100;
    16'b1110111011111100 : data_out = 24'b000000000000000001110100;
    16'b1110111011111101 : data_out = 24'b000000000000000001110100;
    16'b1110111011111110 : data_out = 24'b000000000000000001110100;
    16'b1110111011111111 : data_out = 24'b000000000000000001110100;
    16'b1110111100000000 : data_out = 24'b000000000000000001110100;
    16'b1110111100000001 : data_out = 24'b000000000000000001110100;
    16'b1110111100000010 : data_out = 24'b000000000000000001110101;
    16'b1110111100000011 : data_out = 24'b000000000000000001110101;
    16'b1110111100000100 : data_out = 24'b000000000000000001110101;
    16'b1110111100000101 : data_out = 24'b000000000000000001110101;
    16'b1110111100000110 : data_out = 24'b000000000000000001110101;
    16'b1110111100000111 : data_out = 24'b000000000000000001110101;
    16'b1110111100001000 : data_out = 24'b000000000000000001110101;
    16'b1110111100001001 : data_out = 24'b000000000000000001110101;
    16'b1110111100001010 : data_out = 24'b000000000000000001110101;
    16'b1110111100001011 : data_out = 24'b000000000000000001110110;
    16'b1110111100001100 : data_out = 24'b000000000000000001110110;
    16'b1110111100001101 : data_out = 24'b000000000000000001110110;
    16'b1110111100001110 : data_out = 24'b000000000000000001110110;
    16'b1110111100001111 : data_out = 24'b000000000000000001110110;
    16'b1110111100010000 : data_out = 24'b000000000000000001110110;
    16'b1110111100010001 : data_out = 24'b000000000000000001110110;
    16'b1110111100010010 : data_out = 24'b000000000000000001110110;
    16'b1110111100010011 : data_out = 24'b000000000000000001110111;
    16'b1110111100010100 : data_out = 24'b000000000000000001110111;
    16'b1110111100010101 : data_out = 24'b000000000000000001110111;
    16'b1110111100010110 : data_out = 24'b000000000000000001110111;
    16'b1110111100010111 : data_out = 24'b000000000000000001110111;
    16'b1110111100011000 : data_out = 24'b000000000000000001110111;
    16'b1110111100011001 : data_out = 24'b000000000000000001110111;
    16'b1110111100011010 : data_out = 24'b000000000000000001110111;
    16'b1110111100011011 : data_out = 24'b000000000000000001110111;
    16'b1110111100011100 : data_out = 24'b000000000000000001111000;
    16'b1110111100011101 : data_out = 24'b000000000000000001111000;
    16'b1110111100011110 : data_out = 24'b000000000000000001111000;
    16'b1110111100011111 : data_out = 24'b000000000000000001111000;
    16'b1110111100100000 : data_out = 24'b000000000000000001111000;
    16'b1110111100100001 : data_out = 24'b000000000000000001111000;
    16'b1110111100100010 : data_out = 24'b000000000000000001111000;
    16'b1110111100100011 : data_out = 24'b000000000000000001111000;
    16'b1110111100100100 : data_out = 24'b000000000000000001111001;
    16'b1110111100100101 : data_out = 24'b000000000000000001111001;
    16'b1110111100100110 : data_out = 24'b000000000000000001111001;
    16'b1110111100100111 : data_out = 24'b000000000000000001111001;
    16'b1110111100101000 : data_out = 24'b000000000000000001111001;
    16'b1110111100101001 : data_out = 24'b000000000000000001111001;
    16'b1110111100101010 : data_out = 24'b000000000000000001111001;
    16'b1110111100101011 : data_out = 24'b000000000000000001111001;
    16'b1110111100101100 : data_out = 24'b000000000000000001111001;
    16'b1110111100101101 : data_out = 24'b000000000000000001111010;
    16'b1110111100101110 : data_out = 24'b000000000000000001111010;
    16'b1110111100101111 : data_out = 24'b000000000000000001111010;
    16'b1110111100110000 : data_out = 24'b000000000000000001111010;
    16'b1110111100110001 : data_out = 24'b000000000000000001111010;
    16'b1110111100110010 : data_out = 24'b000000000000000001111010;
    16'b1110111100110011 : data_out = 24'b000000000000000001111010;
    16'b1110111100110100 : data_out = 24'b000000000000000001111010;
    16'b1110111100110101 : data_out = 24'b000000000000000001111011;
    16'b1110111100110110 : data_out = 24'b000000000000000001111011;
    16'b1110111100110111 : data_out = 24'b000000000000000001111011;
    16'b1110111100111000 : data_out = 24'b000000000000000001111011;
    16'b1110111100111001 : data_out = 24'b000000000000000001111011;
    16'b1110111100111010 : data_out = 24'b000000000000000001111011;
    16'b1110111100111011 : data_out = 24'b000000000000000001111011;
    16'b1110111100111100 : data_out = 24'b000000000000000001111011;
    16'b1110111100111101 : data_out = 24'b000000000000000001111100;
    16'b1110111100111110 : data_out = 24'b000000000000000001111100;
    16'b1110111100111111 : data_out = 24'b000000000000000001111100;
    16'b1110111101000000 : data_out = 24'b000000000000000001111100;
    16'b1110111101000001 : data_out = 24'b000000000000000001111100;
    16'b1110111101000010 : data_out = 24'b000000000000000001111100;
    16'b1110111101000011 : data_out = 24'b000000000000000001111100;
    16'b1110111101000100 : data_out = 24'b000000000000000001111100;
    16'b1110111101000101 : data_out = 24'b000000000000000001111100;
    16'b1110111101000110 : data_out = 24'b000000000000000001111101;
    16'b1110111101000111 : data_out = 24'b000000000000000001111101;
    16'b1110111101001000 : data_out = 24'b000000000000000001111101;
    16'b1110111101001001 : data_out = 24'b000000000000000001111101;
    16'b1110111101001010 : data_out = 24'b000000000000000001111101;
    16'b1110111101001011 : data_out = 24'b000000000000000001111101;
    16'b1110111101001100 : data_out = 24'b000000000000000001111101;
    16'b1110111101001101 : data_out = 24'b000000000000000001111101;
    16'b1110111101001110 : data_out = 24'b000000000000000001111110;
    16'b1110111101001111 : data_out = 24'b000000000000000001111110;
    16'b1110111101010000 : data_out = 24'b000000000000000001111110;
    16'b1110111101010001 : data_out = 24'b000000000000000001111110;
    16'b1110111101010010 : data_out = 24'b000000000000000001111110;
    16'b1110111101010011 : data_out = 24'b000000000000000001111110;
    16'b1110111101010100 : data_out = 24'b000000000000000001111110;
    16'b1110111101010101 : data_out = 24'b000000000000000001111110;
    16'b1110111101010110 : data_out = 24'b000000000000000001111111;
    16'b1110111101010111 : data_out = 24'b000000000000000001111111;
    16'b1110111101011000 : data_out = 24'b000000000000000001111111;
    16'b1110111101011001 : data_out = 24'b000000000000000001111111;
    16'b1110111101011010 : data_out = 24'b000000000000000001111111;
    16'b1110111101011011 : data_out = 24'b000000000000000001111111;
    16'b1110111101011100 : data_out = 24'b000000000000000001111111;
    16'b1110111101011101 : data_out = 24'b000000000000000001111111;
    16'b1110111101011110 : data_out = 24'b000000000000000010000000;
    16'b1110111101011111 : data_out = 24'b000000000000000010000000;
    16'b1110111101100000 : data_out = 24'b000000000000000010000000;
    16'b1110111101100001 : data_out = 24'b000000000000000010000000;
    16'b1110111101100010 : data_out = 24'b000000000000000010000000;
    16'b1110111101100011 : data_out = 24'b000000000000000010000000;
    16'b1110111101100100 : data_out = 24'b000000000000000010000000;
    16'b1110111101100101 : data_out = 24'b000000000000000010000000;
    16'b1110111101100110 : data_out = 24'b000000000000000010000001;
    16'b1110111101100111 : data_out = 24'b000000000000000010000001;
    16'b1110111101101000 : data_out = 24'b000000000000000010000001;
    16'b1110111101101001 : data_out = 24'b000000000000000010000001;
    16'b1110111101101010 : data_out = 24'b000000000000000010000001;
    16'b1110111101101011 : data_out = 24'b000000000000000010000001;
    16'b1110111101101100 : data_out = 24'b000000000000000010000001;
    16'b1110111101101101 : data_out = 24'b000000000000000010000001;
    16'b1110111101101110 : data_out = 24'b000000000000000010000010;
    16'b1110111101101111 : data_out = 24'b000000000000000010000010;
    16'b1110111101110000 : data_out = 24'b000000000000000010000010;
    16'b1110111101110001 : data_out = 24'b000000000000000010000010;
    16'b1110111101110010 : data_out = 24'b000000000000000010000010;
    16'b1110111101110011 : data_out = 24'b000000000000000010000010;
    16'b1110111101110100 : data_out = 24'b000000000000000010000010;
    16'b1110111101110101 : data_out = 24'b000000000000000010000010;
    16'b1110111101110110 : data_out = 24'b000000000000000010000011;
    16'b1110111101110111 : data_out = 24'b000000000000000010000011;
    16'b1110111101111000 : data_out = 24'b000000000000000010000011;
    16'b1110111101111001 : data_out = 24'b000000000000000010000011;
    16'b1110111101111010 : data_out = 24'b000000000000000010000011;
    16'b1110111101111011 : data_out = 24'b000000000000000010000011;
    16'b1110111101111100 : data_out = 24'b000000000000000010000011;
    16'b1110111101111101 : data_out = 24'b000000000000000010000100;
    16'b1110111101111110 : data_out = 24'b000000000000000010000100;
    16'b1110111101111111 : data_out = 24'b000000000000000010000100;
    16'b1110111110000000 : data_out = 24'b000000000000000010000100;
    16'b1110111110000001 : data_out = 24'b000000000000000010000100;
    16'b1110111110000010 : data_out = 24'b000000000000000010000100;
    16'b1110111110000011 : data_out = 24'b000000000000000010000100;
    16'b1110111110000100 : data_out = 24'b000000000000000010000100;
    16'b1110111110000101 : data_out = 24'b000000000000000010000101;
    16'b1110111110000110 : data_out = 24'b000000000000000010000101;
    16'b1110111110000111 : data_out = 24'b000000000000000010000101;
    16'b1110111110001000 : data_out = 24'b000000000000000010000101;
    16'b1110111110001001 : data_out = 24'b000000000000000010000101;
    16'b1110111110001010 : data_out = 24'b000000000000000010000101;
    16'b1110111110001011 : data_out = 24'b000000000000000010000101;
    16'b1110111110001100 : data_out = 24'b000000000000000010000101;
    16'b1110111110001101 : data_out = 24'b000000000000000010000110;
    16'b1110111110001110 : data_out = 24'b000000000000000010000110;
    16'b1110111110001111 : data_out = 24'b000000000000000010000110;
    16'b1110111110010000 : data_out = 24'b000000000000000010000110;
    16'b1110111110010001 : data_out = 24'b000000000000000010000110;
    16'b1110111110010010 : data_out = 24'b000000000000000010000110;
    16'b1110111110010011 : data_out = 24'b000000000000000010000110;
    16'b1110111110010100 : data_out = 24'b000000000000000010000111;
    16'b1110111110010101 : data_out = 24'b000000000000000010000111;
    16'b1110111110010110 : data_out = 24'b000000000000000010000111;
    16'b1110111110010111 : data_out = 24'b000000000000000010000111;
    16'b1110111110011000 : data_out = 24'b000000000000000010000111;
    16'b1110111110011001 : data_out = 24'b000000000000000010000111;
    16'b1110111110011010 : data_out = 24'b000000000000000010000111;
    16'b1110111110011011 : data_out = 24'b000000000000000010000111;
    16'b1110111110011100 : data_out = 24'b000000000000000010001000;
    16'b1110111110011101 : data_out = 24'b000000000000000010001000;
    16'b1110111110011110 : data_out = 24'b000000000000000010001000;
    16'b1110111110011111 : data_out = 24'b000000000000000010001000;
    16'b1110111110100000 : data_out = 24'b000000000000000010001000;
    16'b1110111110100001 : data_out = 24'b000000000000000010001000;
    16'b1110111110100010 : data_out = 24'b000000000000000010001000;
    16'b1110111110100011 : data_out = 24'b000000000000000010001001;
    16'b1110111110100100 : data_out = 24'b000000000000000010001001;
    16'b1110111110100101 : data_out = 24'b000000000000000010001001;
    16'b1110111110100110 : data_out = 24'b000000000000000010001001;
    16'b1110111110100111 : data_out = 24'b000000000000000010001001;
    16'b1110111110101000 : data_out = 24'b000000000000000010001001;
    16'b1110111110101001 : data_out = 24'b000000000000000010001001;
    16'b1110111110101010 : data_out = 24'b000000000000000010001001;
    16'b1110111110101011 : data_out = 24'b000000000000000010001010;
    16'b1110111110101100 : data_out = 24'b000000000000000010001010;
    16'b1110111110101101 : data_out = 24'b000000000000000010001010;
    16'b1110111110101110 : data_out = 24'b000000000000000010001010;
    16'b1110111110101111 : data_out = 24'b000000000000000010001010;
    16'b1110111110110000 : data_out = 24'b000000000000000010001010;
    16'b1110111110110001 : data_out = 24'b000000000000000010001010;
    16'b1110111110110010 : data_out = 24'b000000000000000010001011;
    16'b1110111110110011 : data_out = 24'b000000000000000010001011;
    16'b1110111110110100 : data_out = 24'b000000000000000010001011;
    16'b1110111110110101 : data_out = 24'b000000000000000010001011;
    16'b1110111110110110 : data_out = 24'b000000000000000010001011;
    16'b1110111110110111 : data_out = 24'b000000000000000010001011;
    16'b1110111110111000 : data_out = 24'b000000000000000010001011;
    16'b1110111110111001 : data_out = 24'b000000000000000010001011;
    16'b1110111110111010 : data_out = 24'b000000000000000010001100;
    16'b1110111110111011 : data_out = 24'b000000000000000010001100;
    16'b1110111110111100 : data_out = 24'b000000000000000010001100;
    16'b1110111110111101 : data_out = 24'b000000000000000010001100;
    16'b1110111110111110 : data_out = 24'b000000000000000010001100;
    16'b1110111110111111 : data_out = 24'b000000000000000010001100;
    16'b1110111111000000 : data_out = 24'b000000000000000010001100;
    16'b1110111111000001 : data_out = 24'b000000000000000010001101;
    16'b1110111111000010 : data_out = 24'b000000000000000010001101;
    16'b1110111111000011 : data_out = 24'b000000000000000010001101;
    16'b1110111111000100 : data_out = 24'b000000000000000010001101;
    16'b1110111111000101 : data_out = 24'b000000000000000010001101;
    16'b1110111111000110 : data_out = 24'b000000000000000010001101;
    16'b1110111111000111 : data_out = 24'b000000000000000010001101;
    16'b1110111111001000 : data_out = 24'b000000000000000010001110;
    16'b1110111111001001 : data_out = 24'b000000000000000010001110;
    16'b1110111111001010 : data_out = 24'b000000000000000010001110;
    16'b1110111111001011 : data_out = 24'b000000000000000010001110;
    16'b1110111111001100 : data_out = 24'b000000000000000010001110;
    16'b1110111111001101 : data_out = 24'b000000000000000010001110;
    16'b1110111111001110 : data_out = 24'b000000000000000010001110;
    16'b1110111111001111 : data_out = 24'b000000000000000010001111;
    16'b1110111111010000 : data_out = 24'b000000000000000010001111;
    16'b1110111111010001 : data_out = 24'b000000000000000010001111;
    16'b1110111111010010 : data_out = 24'b000000000000000010001111;
    16'b1110111111010011 : data_out = 24'b000000000000000010001111;
    16'b1110111111010100 : data_out = 24'b000000000000000010001111;
    16'b1110111111010101 : data_out = 24'b000000000000000010001111;
    16'b1110111111010110 : data_out = 24'b000000000000000010010000;
    16'b1110111111010111 : data_out = 24'b000000000000000010010000;
    16'b1110111111011000 : data_out = 24'b000000000000000010010000;
    16'b1110111111011001 : data_out = 24'b000000000000000010010000;
    16'b1110111111011010 : data_out = 24'b000000000000000010010000;
    16'b1110111111011011 : data_out = 24'b000000000000000010010000;
    16'b1110111111011100 : data_out = 24'b000000000000000010010000;
    16'b1110111111011101 : data_out = 24'b000000000000000010010000;
    16'b1110111111011110 : data_out = 24'b000000000000000010010001;
    16'b1110111111011111 : data_out = 24'b000000000000000010010001;
    16'b1110111111100000 : data_out = 24'b000000000000000010010001;
    16'b1110111111100001 : data_out = 24'b000000000000000010010001;
    16'b1110111111100010 : data_out = 24'b000000000000000010010001;
    16'b1110111111100011 : data_out = 24'b000000000000000010010001;
    16'b1110111111100100 : data_out = 24'b000000000000000010010001;
    16'b1110111111100101 : data_out = 24'b000000000000000010010010;
    16'b1110111111100110 : data_out = 24'b000000000000000010010010;
    16'b1110111111100111 : data_out = 24'b000000000000000010010010;
    16'b1110111111101000 : data_out = 24'b000000000000000010010010;
    16'b1110111111101001 : data_out = 24'b000000000000000010010010;
    16'b1110111111101010 : data_out = 24'b000000000000000010010010;
    16'b1110111111101011 : data_out = 24'b000000000000000010010010;
    16'b1110111111101100 : data_out = 24'b000000000000000010010011;
    16'b1110111111101101 : data_out = 24'b000000000000000010010011;
    16'b1110111111101110 : data_out = 24'b000000000000000010010011;
    16'b1110111111101111 : data_out = 24'b000000000000000010010011;
    16'b1110111111110000 : data_out = 24'b000000000000000010010011;
    16'b1110111111110001 : data_out = 24'b000000000000000010010011;
    16'b1110111111110010 : data_out = 24'b000000000000000010010100;
    16'b1110111111110011 : data_out = 24'b000000000000000010010100;
    16'b1110111111110100 : data_out = 24'b000000000000000010010100;
    16'b1110111111110101 : data_out = 24'b000000000000000010010100;
    16'b1110111111110110 : data_out = 24'b000000000000000010010100;
    16'b1110111111110111 : data_out = 24'b000000000000000010010100;
    16'b1110111111111000 : data_out = 24'b000000000000000010010100;
    16'b1110111111111001 : data_out = 24'b000000000000000010010101;
    16'b1110111111111010 : data_out = 24'b000000000000000010010101;
    16'b1110111111111011 : data_out = 24'b000000000000000010010101;
    16'b1110111111111100 : data_out = 24'b000000000000000010010101;
    16'b1110111111111101 : data_out = 24'b000000000000000010010101;
    16'b1110111111111110 : data_out = 24'b000000000000000010010101;
    16'b1110111111111111 : data_out = 24'b000000000000000010010101;
    16'b1111000000000000 : data_out = 24'b000000000000000010010110;
    16'b1111000000000001 : data_out = 24'b000000000000000010010110;
    16'b1111000000000010 : data_out = 24'b000000000000000010010110;
    16'b1111000000000011 : data_out = 24'b000000000000000010010110;
    16'b1111000000000100 : data_out = 24'b000000000000000010010110;
    16'b1111000000000101 : data_out = 24'b000000000000000010010110;
    16'b1111000000000110 : data_out = 24'b000000000000000010010110;
    16'b1111000000000111 : data_out = 24'b000000000000000010010111;
    16'b1111000000001000 : data_out = 24'b000000000000000010010111;
    16'b1111000000001001 : data_out = 24'b000000000000000010010111;
    16'b1111000000001010 : data_out = 24'b000000000000000010010111;
    16'b1111000000001011 : data_out = 24'b000000000000000010010111;
    16'b1111000000001100 : data_out = 24'b000000000000000010010111;
    16'b1111000000001101 : data_out = 24'b000000000000000010010111;
    16'b1111000000001110 : data_out = 24'b000000000000000010011000;
    16'b1111000000001111 : data_out = 24'b000000000000000010011000;
    16'b1111000000010000 : data_out = 24'b000000000000000010011000;
    16'b1111000000010001 : data_out = 24'b000000000000000010011000;
    16'b1111000000010010 : data_out = 24'b000000000000000010011000;
    16'b1111000000010011 : data_out = 24'b000000000000000010011000;
    16'b1111000000010100 : data_out = 24'b000000000000000010011001;
    16'b1111000000010101 : data_out = 24'b000000000000000010011001;
    16'b1111000000010110 : data_out = 24'b000000000000000010011001;
    16'b1111000000010111 : data_out = 24'b000000000000000010011001;
    16'b1111000000011000 : data_out = 24'b000000000000000010011001;
    16'b1111000000011001 : data_out = 24'b000000000000000010011001;
    16'b1111000000011010 : data_out = 24'b000000000000000010011001;
    16'b1111000000011011 : data_out = 24'b000000000000000010011010;
    16'b1111000000011100 : data_out = 24'b000000000000000010011010;
    16'b1111000000011101 : data_out = 24'b000000000000000010011010;
    16'b1111000000011110 : data_out = 24'b000000000000000010011010;
    16'b1111000000011111 : data_out = 24'b000000000000000010011010;
    16'b1111000000100000 : data_out = 24'b000000000000000010011010;
    16'b1111000000100001 : data_out = 24'b000000000000000010011010;
    16'b1111000000100010 : data_out = 24'b000000000000000010011011;
    16'b1111000000100011 : data_out = 24'b000000000000000010011011;
    16'b1111000000100100 : data_out = 24'b000000000000000010011011;
    16'b1111000000100101 : data_out = 24'b000000000000000010011011;
    16'b1111000000100110 : data_out = 24'b000000000000000010011011;
    16'b1111000000100111 : data_out = 24'b000000000000000010011011;
    16'b1111000000101000 : data_out = 24'b000000000000000010011100;
    16'b1111000000101001 : data_out = 24'b000000000000000010011100;
    16'b1111000000101010 : data_out = 24'b000000000000000010011100;
    16'b1111000000101011 : data_out = 24'b000000000000000010011100;
    16'b1111000000101100 : data_out = 24'b000000000000000010011100;
    16'b1111000000101101 : data_out = 24'b000000000000000010011100;
    16'b1111000000101110 : data_out = 24'b000000000000000010011100;
    16'b1111000000101111 : data_out = 24'b000000000000000010011101;
    16'b1111000000110000 : data_out = 24'b000000000000000010011101;
    16'b1111000000110001 : data_out = 24'b000000000000000010011101;
    16'b1111000000110010 : data_out = 24'b000000000000000010011101;
    16'b1111000000110011 : data_out = 24'b000000000000000010011101;
    16'b1111000000110100 : data_out = 24'b000000000000000010011101;
    16'b1111000000110101 : data_out = 24'b000000000000000010011110;
    16'b1111000000110110 : data_out = 24'b000000000000000010011110;
    16'b1111000000110111 : data_out = 24'b000000000000000010011110;
    16'b1111000000111000 : data_out = 24'b000000000000000010011110;
    16'b1111000000111001 : data_out = 24'b000000000000000010011110;
    16'b1111000000111010 : data_out = 24'b000000000000000010011110;
    16'b1111000000111011 : data_out = 24'b000000000000000010011110;
    16'b1111000000111100 : data_out = 24'b000000000000000010011111;
    16'b1111000000111101 : data_out = 24'b000000000000000010011111;
    16'b1111000000111110 : data_out = 24'b000000000000000010011111;
    16'b1111000000111111 : data_out = 24'b000000000000000010011111;
    16'b1111000001000000 : data_out = 24'b000000000000000010011111;
    16'b1111000001000001 : data_out = 24'b000000000000000010011111;
    16'b1111000001000010 : data_out = 24'b000000000000000010100000;
    16'b1111000001000011 : data_out = 24'b000000000000000010100000;
    16'b1111000001000100 : data_out = 24'b000000000000000010100000;
    16'b1111000001000101 : data_out = 24'b000000000000000010100000;
    16'b1111000001000110 : data_out = 24'b000000000000000010100000;
    16'b1111000001000111 : data_out = 24'b000000000000000010100000;
    16'b1111000001001000 : data_out = 24'b000000000000000010100000;
    16'b1111000001001001 : data_out = 24'b000000000000000010100001;
    16'b1111000001001010 : data_out = 24'b000000000000000010100001;
    16'b1111000001001011 : data_out = 24'b000000000000000010100001;
    16'b1111000001001100 : data_out = 24'b000000000000000010100001;
    16'b1111000001001101 : data_out = 24'b000000000000000010100001;
    16'b1111000001001110 : data_out = 24'b000000000000000010100001;
    16'b1111000001001111 : data_out = 24'b000000000000000010100010;
    16'b1111000001010000 : data_out = 24'b000000000000000010100010;
    16'b1111000001010001 : data_out = 24'b000000000000000010100010;
    16'b1111000001010010 : data_out = 24'b000000000000000010100010;
    16'b1111000001010011 : data_out = 24'b000000000000000010100010;
    16'b1111000001010100 : data_out = 24'b000000000000000010100010;
    16'b1111000001010101 : data_out = 24'b000000000000000010100011;
    16'b1111000001010110 : data_out = 24'b000000000000000010100011;
    16'b1111000001010111 : data_out = 24'b000000000000000010100011;
    16'b1111000001011000 : data_out = 24'b000000000000000010100011;
    16'b1111000001011001 : data_out = 24'b000000000000000010100011;
    16'b1111000001011010 : data_out = 24'b000000000000000010100011;
    16'b1111000001011011 : data_out = 24'b000000000000000010100011;
    16'b1111000001011100 : data_out = 24'b000000000000000010100100;
    16'b1111000001011101 : data_out = 24'b000000000000000010100100;
    16'b1111000001011110 : data_out = 24'b000000000000000010100100;
    16'b1111000001011111 : data_out = 24'b000000000000000010100100;
    16'b1111000001100000 : data_out = 24'b000000000000000010100100;
    16'b1111000001100001 : data_out = 24'b000000000000000010100100;
    16'b1111000001100010 : data_out = 24'b000000000000000010100101;
    16'b1111000001100011 : data_out = 24'b000000000000000010100101;
    16'b1111000001100100 : data_out = 24'b000000000000000010100101;
    16'b1111000001100101 : data_out = 24'b000000000000000010100101;
    16'b1111000001100110 : data_out = 24'b000000000000000010100101;
    16'b1111000001100111 : data_out = 24'b000000000000000010100101;
    16'b1111000001101000 : data_out = 24'b000000000000000010100110;
    16'b1111000001101001 : data_out = 24'b000000000000000010100110;
    16'b1111000001101010 : data_out = 24'b000000000000000010100110;
    16'b1111000001101011 : data_out = 24'b000000000000000010100110;
    16'b1111000001101100 : data_out = 24'b000000000000000010100110;
    16'b1111000001101101 : data_out = 24'b000000000000000010100110;
    16'b1111000001101110 : data_out = 24'b000000000000000010100111;
    16'b1111000001101111 : data_out = 24'b000000000000000010100111;
    16'b1111000001110000 : data_out = 24'b000000000000000010100111;
    16'b1111000001110001 : data_out = 24'b000000000000000010100111;
    16'b1111000001110010 : data_out = 24'b000000000000000010100111;
    16'b1111000001110011 : data_out = 24'b000000000000000010100111;
    16'b1111000001110100 : data_out = 24'b000000000000000010101000;
    16'b1111000001110101 : data_out = 24'b000000000000000010101000;
    16'b1111000001110110 : data_out = 24'b000000000000000010101000;
    16'b1111000001110111 : data_out = 24'b000000000000000010101000;
    16'b1111000001111000 : data_out = 24'b000000000000000010101000;
    16'b1111000001111001 : data_out = 24'b000000000000000010101000;
    16'b1111000001111010 : data_out = 24'b000000000000000010101001;
    16'b1111000001111011 : data_out = 24'b000000000000000010101001;
    16'b1111000001111100 : data_out = 24'b000000000000000010101001;
    16'b1111000001111101 : data_out = 24'b000000000000000010101001;
    16'b1111000001111110 : data_out = 24'b000000000000000010101001;
    16'b1111000001111111 : data_out = 24'b000000000000000010101001;
    16'b1111000010000000 : data_out = 24'b000000000000000010101010;
    16'b1111000010000001 : data_out = 24'b000000000000000010101010;
    16'b1111000010000010 : data_out = 24'b000000000000000010101010;
    16'b1111000010000011 : data_out = 24'b000000000000000010101010;
    16'b1111000010000100 : data_out = 24'b000000000000000010101010;
    16'b1111000010000101 : data_out = 24'b000000000000000010101010;
    16'b1111000010000110 : data_out = 24'b000000000000000010101011;
    16'b1111000010000111 : data_out = 24'b000000000000000010101011;
    16'b1111000010001000 : data_out = 24'b000000000000000010101011;
    16'b1111000010001001 : data_out = 24'b000000000000000010101011;
    16'b1111000010001010 : data_out = 24'b000000000000000010101011;
    16'b1111000010001011 : data_out = 24'b000000000000000010101011;
    16'b1111000010001100 : data_out = 24'b000000000000000010101100;
    16'b1111000010001101 : data_out = 24'b000000000000000010101100;
    16'b1111000010001110 : data_out = 24'b000000000000000010101100;
    16'b1111000010001111 : data_out = 24'b000000000000000010101100;
    16'b1111000010010000 : data_out = 24'b000000000000000010101100;
    16'b1111000010010001 : data_out = 24'b000000000000000010101100;
    16'b1111000010010010 : data_out = 24'b000000000000000010101101;
    16'b1111000010010011 : data_out = 24'b000000000000000010101101;
    16'b1111000010010100 : data_out = 24'b000000000000000010101101;
    16'b1111000010010101 : data_out = 24'b000000000000000010101101;
    16'b1111000010010110 : data_out = 24'b000000000000000010101101;
    16'b1111000010010111 : data_out = 24'b000000000000000010101101;
    16'b1111000010011000 : data_out = 24'b000000000000000010101110;
    16'b1111000010011001 : data_out = 24'b000000000000000010101110;
    16'b1111000010011010 : data_out = 24'b000000000000000010101110;
    16'b1111000010011011 : data_out = 24'b000000000000000010101110;
    16'b1111000010011100 : data_out = 24'b000000000000000010101110;
    16'b1111000010011101 : data_out = 24'b000000000000000010101110;
    16'b1111000010011110 : data_out = 24'b000000000000000010101111;
    16'b1111000010011111 : data_out = 24'b000000000000000010101111;
    16'b1111000010100000 : data_out = 24'b000000000000000010101111;
    16'b1111000010100001 : data_out = 24'b000000000000000010101111;
    16'b1111000010100010 : data_out = 24'b000000000000000010101111;
    16'b1111000010100011 : data_out = 24'b000000000000000010101111;
    16'b1111000010100100 : data_out = 24'b000000000000000010110000;
    16'b1111000010100101 : data_out = 24'b000000000000000010110000;
    16'b1111000010100110 : data_out = 24'b000000000000000010110000;
    16'b1111000010100111 : data_out = 24'b000000000000000010110000;
    16'b1111000010101000 : data_out = 24'b000000000000000010110000;
    16'b1111000010101001 : data_out = 24'b000000000000000010110000;
    16'b1111000010101010 : data_out = 24'b000000000000000010110001;
    16'b1111000010101011 : data_out = 24'b000000000000000010110001;
    16'b1111000010101100 : data_out = 24'b000000000000000010110001;
    16'b1111000010101101 : data_out = 24'b000000000000000010110001;
    16'b1111000010101110 : data_out = 24'b000000000000000010110001;
    16'b1111000010101111 : data_out = 24'b000000000000000010110010;
    16'b1111000010110000 : data_out = 24'b000000000000000010110010;
    16'b1111000010110001 : data_out = 24'b000000000000000010110010;
    16'b1111000010110010 : data_out = 24'b000000000000000010110010;
    16'b1111000010110011 : data_out = 24'b000000000000000010110010;
    16'b1111000010110100 : data_out = 24'b000000000000000010110010;
    16'b1111000010110101 : data_out = 24'b000000000000000010110011;
    16'b1111000010110110 : data_out = 24'b000000000000000010110011;
    16'b1111000010110111 : data_out = 24'b000000000000000010110011;
    16'b1111000010111000 : data_out = 24'b000000000000000010110011;
    16'b1111000010111001 : data_out = 24'b000000000000000010110011;
    16'b1111000010111010 : data_out = 24'b000000000000000010110011;
    16'b1111000010111011 : data_out = 24'b000000000000000010110100;
    16'b1111000010111100 : data_out = 24'b000000000000000010110100;
    16'b1111000010111101 : data_out = 24'b000000000000000010110100;
    16'b1111000010111110 : data_out = 24'b000000000000000010110100;
    16'b1111000010111111 : data_out = 24'b000000000000000010110100;
    16'b1111000011000000 : data_out = 24'b000000000000000010110100;
    16'b1111000011000001 : data_out = 24'b000000000000000010110101;
    16'b1111000011000010 : data_out = 24'b000000000000000010110101;
    16'b1111000011000011 : data_out = 24'b000000000000000010110101;
    16'b1111000011000100 : data_out = 24'b000000000000000010110101;
    16'b1111000011000101 : data_out = 24'b000000000000000010110101;
    16'b1111000011000110 : data_out = 24'b000000000000000010110110;
    16'b1111000011000111 : data_out = 24'b000000000000000010110110;
    16'b1111000011001000 : data_out = 24'b000000000000000010110110;
    16'b1111000011001001 : data_out = 24'b000000000000000010110110;
    16'b1111000011001010 : data_out = 24'b000000000000000010110110;
    16'b1111000011001011 : data_out = 24'b000000000000000010110110;
    16'b1111000011001100 : data_out = 24'b000000000000000010110111;
    16'b1111000011001101 : data_out = 24'b000000000000000010110111;
    16'b1111000011001110 : data_out = 24'b000000000000000010110111;
    16'b1111000011001111 : data_out = 24'b000000000000000010110111;
    16'b1111000011010000 : data_out = 24'b000000000000000010110111;
    16'b1111000011010001 : data_out = 24'b000000000000000010111000;
    16'b1111000011010010 : data_out = 24'b000000000000000010111000;
    16'b1111000011010011 : data_out = 24'b000000000000000010111000;
    16'b1111000011010100 : data_out = 24'b000000000000000010111000;
    16'b1111000011010101 : data_out = 24'b000000000000000010111000;
    16'b1111000011010110 : data_out = 24'b000000000000000010111000;
    16'b1111000011010111 : data_out = 24'b000000000000000010111001;
    16'b1111000011011000 : data_out = 24'b000000000000000010111001;
    16'b1111000011011001 : data_out = 24'b000000000000000010111001;
    16'b1111000011011010 : data_out = 24'b000000000000000010111001;
    16'b1111000011011011 : data_out = 24'b000000000000000010111001;
    16'b1111000011011100 : data_out = 24'b000000000000000010111010;
    16'b1111000011011101 : data_out = 24'b000000000000000010111010;
    16'b1111000011011110 : data_out = 24'b000000000000000010111010;
    16'b1111000011011111 : data_out = 24'b000000000000000010111010;
    16'b1111000011100000 : data_out = 24'b000000000000000010111010;
    16'b1111000011100001 : data_out = 24'b000000000000000010111010;
    16'b1111000011100010 : data_out = 24'b000000000000000010111011;
    16'b1111000011100011 : data_out = 24'b000000000000000010111011;
    16'b1111000011100100 : data_out = 24'b000000000000000010111011;
    16'b1111000011100101 : data_out = 24'b000000000000000010111011;
    16'b1111000011100110 : data_out = 24'b000000000000000010111011;
    16'b1111000011100111 : data_out = 24'b000000000000000010111100;
    16'b1111000011101000 : data_out = 24'b000000000000000010111100;
    16'b1111000011101001 : data_out = 24'b000000000000000010111100;
    16'b1111000011101010 : data_out = 24'b000000000000000010111100;
    16'b1111000011101011 : data_out = 24'b000000000000000010111100;
    16'b1111000011101100 : data_out = 24'b000000000000000010111100;
    16'b1111000011101101 : data_out = 24'b000000000000000010111101;
    16'b1111000011101110 : data_out = 24'b000000000000000010111101;
    16'b1111000011101111 : data_out = 24'b000000000000000010111101;
    16'b1111000011110000 : data_out = 24'b000000000000000010111101;
    16'b1111000011110001 : data_out = 24'b000000000000000010111101;
    16'b1111000011110010 : data_out = 24'b000000000000000010111110;
    16'b1111000011110011 : data_out = 24'b000000000000000010111110;
    16'b1111000011110100 : data_out = 24'b000000000000000010111110;
    16'b1111000011110101 : data_out = 24'b000000000000000010111110;
    16'b1111000011110110 : data_out = 24'b000000000000000010111110;
    16'b1111000011110111 : data_out = 24'b000000000000000010111110;
    16'b1111000011111000 : data_out = 24'b000000000000000010111111;
    16'b1111000011111001 : data_out = 24'b000000000000000010111111;
    16'b1111000011111010 : data_out = 24'b000000000000000010111111;
    16'b1111000011111011 : data_out = 24'b000000000000000010111111;
    16'b1111000011111100 : data_out = 24'b000000000000000010111111;
    16'b1111000011111101 : data_out = 24'b000000000000000011000000;
    16'b1111000011111110 : data_out = 24'b000000000000000011000000;
    16'b1111000011111111 : data_out = 24'b000000000000000011000000;
    16'b1111000100000000 : data_out = 24'b000000000000000011000000;
    16'b1111000100000001 : data_out = 24'b000000000000000011000000;
    16'b1111000100000010 : data_out = 24'b000000000000000011000001;
    16'b1111000100000011 : data_out = 24'b000000000000000011000001;
    16'b1111000100000100 : data_out = 24'b000000000000000011000001;
    16'b1111000100000101 : data_out = 24'b000000000000000011000001;
    16'b1111000100000110 : data_out = 24'b000000000000000011000001;
    16'b1111000100000111 : data_out = 24'b000000000000000011000001;
    16'b1111000100001000 : data_out = 24'b000000000000000011000010;
    16'b1111000100001001 : data_out = 24'b000000000000000011000010;
    16'b1111000100001010 : data_out = 24'b000000000000000011000010;
    16'b1111000100001011 : data_out = 24'b000000000000000011000010;
    16'b1111000100001100 : data_out = 24'b000000000000000011000010;
    16'b1111000100001101 : data_out = 24'b000000000000000011000011;
    16'b1111000100001110 : data_out = 24'b000000000000000011000011;
    16'b1111000100001111 : data_out = 24'b000000000000000011000011;
    16'b1111000100010000 : data_out = 24'b000000000000000011000011;
    16'b1111000100010001 : data_out = 24'b000000000000000011000011;
    16'b1111000100010010 : data_out = 24'b000000000000000011000100;
    16'b1111000100010011 : data_out = 24'b000000000000000011000100;
    16'b1111000100010100 : data_out = 24'b000000000000000011000100;
    16'b1111000100010101 : data_out = 24'b000000000000000011000100;
    16'b1111000100010110 : data_out = 24'b000000000000000011000100;
    16'b1111000100010111 : data_out = 24'b000000000000000011000101;
    16'b1111000100011000 : data_out = 24'b000000000000000011000101;
    16'b1111000100011001 : data_out = 24'b000000000000000011000101;
    16'b1111000100011010 : data_out = 24'b000000000000000011000101;
    16'b1111000100011011 : data_out = 24'b000000000000000011000101;
    16'b1111000100011100 : data_out = 24'b000000000000000011000101;
    16'b1111000100011101 : data_out = 24'b000000000000000011000110;
    16'b1111000100011110 : data_out = 24'b000000000000000011000110;
    16'b1111000100011111 : data_out = 24'b000000000000000011000110;
    16'b1111000100100000 : data_out = 24'b000000000000000011000110;
    16'b1111000100100001 : data_out = 24'b000000000000000011000110;
    16'b1111000100100010 : data_out = 24'b000000000000000011000111;
    16'b1111000100100011 : data_out = 24'b000000000000000011000111;
    16'b1111000100100100 : data_out = 24'b000000000000000011000111;
    16'b1111000100100101 : data_out = 24'b000000000000000011000111;
    16'b1111000100100110 : data_out = 24'b000000000000000011000111;
    16'b1111000100100111 : data_out = 24'b000000000000000011001000;
    16'b1111000100101000 : data_out = 24'b000000000000000011001000;
    16'b1111000100101001 : data_out = 24'b000000000000000011001000;
    16'b1111000100101010 : data_out = 24'b000000000000000011001000;
    16'b1111000100101011 : data_out = 24'b000000000000000011001000;
    16'b1111000100101100 : data_out = 24'b000000000000000011001001;
    16'b1111000100101101 : data_out = 24'b000000000000000011001001;
    16'b1111000100101110 : data_out = 24'b000000000000000011001001;
    16'b1111000100101111 : data_out = 24'b000000000000000011001001;
    16'b1111000100110000 : data_out = 24'b000000000000000011001001;
    16'b1111000100110001 : data_out = 24'b000000000000000011001010;
    16'b1111000100110010 : data_out = 24'b000000000000000011001010;
    16'b1111000100110011 : data_out = 24'b000000000000000011001010;
    16'b1111000100110100 : data_out = 24'b000000000000000011001010;
    16'b1111000100110101 : data_out = 24'b000000000000000011001010;
    16'b1111000100110110 : data_out = 24'b000000000000000011001011;
    16'b1111000100110111 : data_out = 24'b000000000000000011001011;
    16'b1111000100111000 : data_out = 24'b000000000000000011001011;
    16'b1111000100111001 : data_out = 24'b000000000000000011001011;
    16'b1111000100111010 : data_out = 24'b000000000000000011001011;
    16'b1111000100111011 : data_out = 24'b000000000000000011001100;
    16'b1111000100111100 : data_out = 24'b000000000000000011001100;
    16'b1111000100111101 : data_out = 24'b000000000000000011001100;
    16'b1111000100111110 : data_out = 24'b000000000000000011001100;
    16'b1111000100111111 : data_out = 24'b000000000000000011001100;
    16'b1111000101000000 : data_out = 24'b000000000000000011001101;
    16'b1111000101000001 : data_out = 24'b000000000000000011001101;
    16'b1111000101000010 : data_out = 24'b000000000000000011001101;
    16'b1111000101000011 : data_out = 24'b000000000000000011001101;
    16'b1111000101000100 : data_out = 24'b000000000000000011001101;
    16'b1111000101000101 : data_out = 24'b000000000000000011001110;
    16'b1111000101000110 : data_out = 24'b000000000000000011001110;
    16'b1111000101000111 : data_out = 24'b000000000000000011001110;
    16'b1111000101001000 : data_out = 24'b000000000000000011001110;
    16'b1111000101001001 : data_out = 24'b000000000000000011001110;
    16'b1111000101001010 : data_out = 24'b000000000000000011001111;
    16'b1111000101001011 : data_out = 24'b000000000000000011001111;
    16'b1111000101001100 : data_out = 24'b000000000000000011001111;
    16'b1111000101001101 : data_out = 24'b000000000000000011001111;
    16'b1111000101001110 : data_out = 24'b000000000000000011001111;
    16'b1111000101001111 : data_out = 24'b000000000000000011010000;
    16'b1111000101010000 : data_out = 24'b000000000000000011010000;
    16'b1111000101010001 : data_out = 24'b000000000000000011010000;
    16'b1111000101010010 : data_out = 24'b000000000000000011010000;
    16'b1111000101010011 : data_out = 24'b000000000000000011010000;
    16'b1111000101010100 : data_out = 24'b000000000000000011010001;
    16'b1111000101010101 : data_out = 24'b000000000000000011010001;
    16'b1111000101010110 : data_out = 24'b000000000000000011010001;
    16'b1111000101010111 : data_out = 24'b000000000000000011010001;
    16'b1111000101011000 : data_out = 24'b000000000000000011010001;
    16'b1111000101011001 : data_out = 24'b000000000000000011010010;
    16'b1111000101011010 : data_out = 24'b000000000000000011010010;
    16'b1111000101011011 : data_out = 24'b000000000000000011010010;
    16'b1111000101011100 : data_out = 24'b000000000000000011010010;
    16'b1111000101011101 : data_out = 24'b000000000000000011010010;
    16'b1111000101011110 : data_out = 24'b000000000000000011010011;
    16'b1111000101011111 : data_out = 24'b000000000000000011010011;
    16'b1111000101100000 : data_out = 24'b000000000000000011010011;
    16'b1111000101100001 : data_out = 24'b000000000000000011010011;
    16'b1111000101100010 : data_out = 24'b000000000000000011010100;
    16'b1111000101100011 : data_out = 24'b000000000000000011010100;
    16'b1111000101100100 : data_out = 24'b000000000000000011010100;
    16'b1111000101100101 : data_out = 24'b000000000000000011010100;
    16'b1111000101100110 : data_out = 24'b000000000000000011010100;
    16'b1111000101100111 : data_out = 24'b000000000000000011010101;
    16'b1111000101101000 : data_out = 24'b000000000000000011010101;
    16'b1111000101101001 : data_out = 24'b000000000000000011010101;
    16'b1111000101101010 : data_out = 24'b000000000000000011010101;
    16'b1111000101101011 : data_out = 24'b000000000000000011010101;
    16'b1111000101101100 : data_out = 24'b000000000000000011010110;
    16'b1111000101101101 : data_out = 24'b000000000000000011010110;
    16'b1111000101101110 : data_out = 24'b000000000000000011010110;
    16'b1111000101101111 : data_out = 24'b000000000000000011010110;
    16'b1111000101110000 : data_out = 24'b000000000000000011010110;
    16'b1111000101110001 : data_out = 24'b000000000000000011010111;
    16'b1111000101110010 : data_out = 24'b000000000000000011010111;
    16'b1111000101110011 : data_out = 24'b000000000000000011010111;
    16'b1111000101110100 : data_out = 24'b000000000000000011010111;
    16'b1111000101110101 : data_out = 24'b000000000000000011010111;
    16'b1111000101110110 : data_out = 24'b000000000000000011011000;
    16'b1111000101110111 : data_out = 24'b000000000000000011011000;
    16'b1111000101111000 : data_out = 24'b000000000000000011011000;
    16'b1111000101111001 : data_out = 24'b000000000000000011011000;
    16'b1111000101111010 : data_out = 24'b000000000000000011011001;
    16'b1111000101111011 : data_out = 24'b000000000000000011011001;
    16'b1111000101111100 : data_out = 24'b000000000000000011011001;
    16'b1111000101111101 : data_out = 24'b000000000000000011011001;
    16'b1111000101111110 : data_out = 24'b000000000000000011011001;
    16'b1111000101111111 : data_out = 24'b000000000000000011011010;
    16'b1111000110000000 : data_out = 24'b000000000000000011011010;
    16'b1111000110000001 : data_out = 24'b000000000000000011011010;
    16'b1111000110000010 : data_out = 24'b000000000000000011011010;
    16'b1111000110000011 : data_out = 24'b000000000000000011011010;
    16'b1111000110000100 : data_out = 24'b000000000000000011011011;
    16'b1111000110000101 : data_out = 24'b000000000000000011011011;
    16'b1111000110000110 : data_out = 24'b000000000000000011011011;
    16'b1111000110000111 : data_out = 24'b000000000000000011011011;
    16'b1111000110001000 : data_out = 24'b000000000000000011011100;
    16'b1111000110001001 : data_out = 24'b000000000000000011011100;
    16'b1111000110001010 : data_out = 24'b000000000000000011011100;
    16'b1111000110001011 : data_out = 24'b000000000000000011011100;
    16'b1111000110001100 : data_out = 24'b000000000000000011011100;
    16'b1111000110001101 : data_out = 24'b000000000000000011011101;
    16'b1111000110001110 : data_out = 24'b000000000000000011011101;
    16'b1111000110001111 : data_out = 24'b000000000000000011011101;
    16'b1111000110010000 : data_out = 24'b000000000000000011011101;
    16'b1111000110010001 : data_out = 24'b000000000000000011011101;
    16'b1111000110010010 : data_out = 24'b000000000000000011011110;
    16'b1111000110010011 : data_out = 24'b000000000000000011011110;
    16'b1111000110010100 : data_out = 24'b000000000000000011011110;
    16'b1111000110010101 : data_out = 24'b000000000000000011011110;
    16'b1111000110010110 : data_out = 24'b000000000000000011011111;
    16'b1111000110010111 : data_out = 24'b000000000000000011011111;
    16'b1111000110011000 : data_out = 24'b000000000000000011011111;
    16'b1111000110011001 : data_out = 24'b000000000000000011011111;
    16'b1111000110011010 : data_out = 24'b000000000000000011011111;
    16'b1111000110011011 : data_out = 24'b000000000000000011100000;
    16'b1111000110011100 : data_out = 24'b000000000000000011100000;
    16'b1111000110011101 : data_out = 24'b000000000000000011100000;
    16'b1111000110011110 : data_out = 24'b000000000000000011100000;
    16'b1111000110011111 : data_out = 24'b000000000000000011100001;
    16'b1111000110100000 : data_out = 24'b000000000000000011100001;
    16'b1111000110100001 : data_out = 24'b000000000000000011100001;
    16'b1111000110100010 : data_out = 24'b000000000000000011100001;
    16'b1111000110100011 : data_out = 24'b000000000000000011100001;
    16'b1111000110100100 : data_out = 24'b000000000000000011100010;
    16'b1111000110100101 : data_out = 24'b000000000000000011100010;
    16'b1111000110100110 : data_out = 24'b000000000000000011100010;
    16'b1111000110100111 : data_out = 24'b000000000000000011100010;
    16'b1111000110101000 : data_out = 24'b000000000000000011100011;
    16'b1111000110101001 : data_out = 24'b000000000000000011100011;
    16'b1111000110101010 : data_out = 24'b000000000000000011100011;
    16'b1111000110101011 : data_out = 24'b000000000000000011100011;
    16'b1111000110101100 : data_out = 24'b000000000000000011100011;
    16'b1111000110101101 : data_out = 24'b000000000000000011100100;
    16'b1111000110101110 : data_out = 24'b000000000000000011100100;
    16'b1111000110101111 : data_out = 24'b000000000000000011100100;
    16'b1111000110110000 : data_out = 24'b000000000000000011100100;
    16'b1111000110110001 : data_out = 24'b000000000000000011100101;
    16'b1111000110110010 : data_out = 24'b000000000000000011100101;
    16'b1111000110110011 : data_out = 24'b000000000000000011100101;
    16'b1111000110110100 : data_out = 24'b000000000000000011100101;
    16'b1111000110110101 : data_out = 24'b000000000000000011100101;
    16'b1111000110110110 : data_out = 24'b000000000000000011100110;
    16'b1111000110110111 : data_out = 24'b000000000000000011100110;
    16'b1111000110111000 : data_out = 24'b000000000000000011100110;
    16'b1111000110111001 : data_out = 24'b000000000000000011100110;
    16'b1111000110111010 : data_out = 24'b000000000000000011100111;
    16'b1111000110111011 : data_out = 24'b000000000000000011100111;
    16'b1111000110111100 : data_out = 24'b000000000000000011100111;
    16'b1111000110111101 : data_out = 24'b000000000000000011100111;
    16'b1111000110111110 : data_out = 24'b000000000000000011100111;
    16'b1111000110111111 : data_out = 24'b000000000000000011101000;
    16'b1111000111000000 : data_out = 24'b000000000000000011101000;
    16'b1111000111000001 : data_out = 24'b000000000000000011101000;
    16'b1111000111000010 : data_out = 24'b000000000000000011101000;
    16'b1111000111000011 : data_out = 24'b000000000000000011101001;
    16'b1111000111000100 : data_out = 24'b000000000000000011101001;
    16'b1111000111000101 : data_out = 24'b000000000000000011101001;
    16'b1111000111000110 : data_out = 24'b000000000000000011101001;
    16'b1111000111000111 : data_out = 24'b000000000000000011101001;
    16'b1111000111001000 : data_out = 24'b000000000000000011101010;
    16'b1111000111001001 : data_out = 24'b000000000000000011101010;
    16'b1111000111001010 : data_out = 24'b000000000000000011101010;
    16'b1111000111001011 : data_out = 24'b000000000000000011101010;
    16'b1111000111001100 : data_out = 24'b000000000000000011101011;
    16'b1111000111001101 : data_out = 24'b000000000000000011101011;
    16'b1111000111001110 : data_out = 24'b000000000000000011101011;
    16'b1111000111001111 : data_out = 24'b000000000000000011101011;
    16'b1111000111010000 : data_out = 24'b000000000000000011101100;
    16'b1111000111010001 : data_out = 24'b000000000000000011101100;
    16'b1111000111010010 : data_out = 24'b000000000000000011101100;
    16'b1111000111010011 : data_out = 24'b000000000000000011101100;
    16'b1111000111010100 : data_out = 24'b000000000000000011101100;
    16'b1111000111010101 : data_out = 24'b000000000000000011101101;
    16'b1111000111010110 : data_out = 24'b000000000000000011101101;
    16'b1111000111010111 : data_out = 24'b000000000000000011101101;
    16'b1111000111011000 : data_out = 24'b000000000000000011101101;
    16'b1111000111011001 : data_out = 24'b000000000000000011101110;
    16'b1111000111011010 : data_out = 24'b000000000000000011101110;
    16'b1111000111011011 : data_out = 24'b000000000000000011101110;
    16'b1111000111011100 : data_out = 24'b000000000000000011101110;
    16'b1111000111011101 : data_out = 24'b000000000000000011101111;
    16'b1111000111011110 : data_out = 24'b000000000000000011101111;
    16'b1111000111011111 : data_out = 24'b000000000000000011101111;
    16'b1111000111100000 : data_out = 24'b000000000000000011101111;
    16'b1111000111100001 : data_out = 24'b000000000000000011110000;
    16'b1111000111100010 : data_out = 24'b000000000000000011110000;
    16'b1111000111100011 : data_out = 24'b000000000000000011110000;
    16'b1111000111100100 : data_out = 24'b000000000000000011110000;
    16'b1111000111100101 : data_out = 24'b000000000000000011110000;
    16'b1111000111100110 : data_out = 24'b000000000000000011110001;
    16'b1111000111100111 : data_out = 24'b000000000000000011110001;
    16'b1111000111101000 : data_out = 24'b000000000000000011110001;
    16'b1111000111101001 : data_out = 24'b000000000000000011110001;
    16'b1111000111101010 : data_out = 24'b000000000000000011110010;
    16'b1111000111101011 : data_out = 24'b000000000000000011110010;
    16'b1111000111101100 : data_out = 24'b000000000000000011110010;
    16'b1111000111101101 : data_out = 24'b000000000000000011110010;
    16'b1111000111101110 : data_out = 24'b000000000000000011110011;
    16'b1111000111101111 : data_out = 24'b000000000000000011110011;
    16'b1111000111110000 : data_out = 24'b000000000000000011110011;
    16'b1111000111110001 : data_out = 24'b000000000000000011110011;
    16'b1111000111110010 : data_out = 24'b000000000000000011110100;
    16'b1111000111110011 : data_out = 24'b000000000000000011110100;
    16'b1111000111110100 : data_out = 24'b000000000000000011110100;
    16'b1111000111110101 : data_out = 24'b000000000000000011110100;
    16'b1111000111110110 : data_out = 24'b000000000000000011110100;
    16'b1111000111110111 : data_out = 24'b000000000000000011110101;
    16'b1111000111111000 : data_out = 24'b000000000000000011110101;
    16'b1111000111111001 : data_out = 24'b000000000000000011110101;
    16'b1111000111111010 : data_out = 24'b000000000000000011110101;
    16'b1111000111111011 : data_out = 24'b000000000000000011110110;
    16'b1111000111111100 : data_out = 24'b000000000000000011110110;
    16'b1111000111111101 : data_out = 24'b000000000000000011110110;
    16'b1111000111111110 : data_out = 24'b000000000000000011110110;
    16'b1111000111111111 : data_out = 24'b000000000000000011110111;
    16'b1111001000000000 : data_out = 24'b000000000000000011110111;
    16'b1111001000000001 : data_out = 24'b000000000000000011110111;
    16'b1111001000000010 : data_out = 24'b000000000000000011110111;
    16'b1111001000000011 : data_out = 24'b000000000000000011111000;
    16'b1111001000000100 : data_out = 24'b000000000000000011111000;
    16'b1111001000000101 : data_out = 24'b000000000000000011111000;
    16'b1111001000000110 : data_out = 24'b000000000000000011111000;
    16'b1111001000000111 : data_out = 24'b000000000000000011111001;
    16'b1111001000001000 : data_out = 24'b000000000000000011111001;
    16'b1111001000001001 : data_out = 24'b000000000000000011111001;
    16'b1111001000001010 : data_out = 24'b000000000000000011111001;
    16'b1111001000001011 : data_out = 24'b000000000000000011111010;
    16'b1111001000001100 : data_out = 24'b000000000000000011111010;
    16'b1111001000001101 : data_out = 24'b000000000000000011111010;
    16'b1111001000001110 : data_out = 24'b000000000000000011111010;
    16'b1111001000001111 : data_out = 24'b000000000000000011111011;
    16'b1111001000010000 : data_out = 24'b000000000000000011111011;
    16'b1111001000010001 : data_out = 24'b000000000000000011111011;
    16'b1111001000010010 : data_out = 24'b000000000000000011111011;
    16'b1111001000010011 : data_out = 24'b000000000000000011111100;
    16'b1111001000010100 : data_out = 24'b000000000000000011111100;
    16'b1111001000010101 : data_out = 24'b000000000000000011111100;
    16'b1111001000010110 : data_out = 24'b000000000000000011111100;
    16'b1111001000010111 : data_out = 24'b000000000000000011111100;
    16'b1111001000011000 : data_out = 24'b000000000000000011111101;
    16'b1111001000011001 : data_out = 24'b000000000000000011111101;
    16'b1111001000011010 : data_out = 24'b000000000000000011111101;
    16'b1111001000011011 : data_out = 24'b000000000000000011111101;
    16'b1111001000011100 : data_out = 24'b000000000000000011111110;
    16'b1111001000011101 : data_out = 24'b000000000000000011111110;
    16'b1111001000011110 : data_out = 24'b000000000000000011111110;
    16'b1111001000011111 : data_out = 24'b000000000000000011111110;
    16'b1111001000100000 : data_out = 24'b000000000000000011111111;
    16'b1111001000100001 : data_out = 24'b000000000000000011111111;
    16'b1111001000100010 : data_out = 24'b000000000000000011111111;
    16'b1111001000100011 : data_out = 24'b000000000000000011111111;
    16'b1111001000100100 : data_out = 24'b000000000000000100000000;
    16'b1111001000100101 : data_out = 24'b000000000000000100000000;
    16'b1111001000100110 : data_out = 24'b000000000000000100000000;
    16'b1111001000100111 : data_out = 24'b000000000000000100000000;
    16'b1111001000101000 : data_out = 24'b000000000000000100000001;
    16'b1111001000101001 : data_out = 24'b000000000000000100000001;
    16'b1111001000101010 : data_out = 24'b000000000000000100000001;
    16'b1111001000101011 : data_out = 24'b000000000000000100000001;
    16'b1111001000101100 : data_out = 24'b000000000000000100000010;
    16'b1111001000101101 : data_out = 24'b000000000000000100000010;
    16'b1111001000101110 : data_out = 24'b000000000000000100000010;
    16'b1111001000101111 : data_out = 24'b000000000000000100000010;
    16'b1111001000110000 : data_out = 24'b000000000000000100000011;
    16'b1111001000110001 : data_out = 24'b000000000000000100000011;
    16'b1111001000110010 : data_out = 24'b000000000000000100000011;
    16'b1111001000110011 : data_out = 24'b000000000000000100000100;
    16'b1111001000110100 : data_out = 24'b000000000000000100000100;
    16'b1111001000110101 : data_out = 24'b000000000000000100000100;
    16'b1111001000110110 : data_out = 24'b000000000000000100000100;
    16'b1111001000110111 : data_out = 24'b000000000000000100000101;
    16'b1111001000111000 : data_out = 24'b000000000000000100000101;
    16'b1111001000111001 : data_out = 24'b000000000000000100000101;
    16'b1111001000111010 : data_out = 24'b000000000000000100000101;
    16'b1111001000111011 : data_out = 24'b000000000000000100000110;
    16'b1111001000111100 : data_out = 24'b000000000000000100000110;
    16'b1111001000111101 : data_out = 24'b000000000000000100000110;
    16'b1111001000111110 : data_out = 24'b000000000000000100000110;
    16'b1111001000111111 : data_out = 24'b000000000000000100000111;
    16'b1111001001000000 : data_out = 24'b000000000000000100000111;
    16'b1111001001000001 : data_out = 24'b000000000000000100000111;
    16'b1111001001000010 : data_out = 24'b000000000000000100000111;
    16'b1111001001000011 : data_out = 24'b000000000000000100001000;
    16'b1111001001000100 : data_out = 24'b000000000000000100001000;
    16'b1111001001000101 : data_out = 24'b000000000000000100001000;
    16'b1111001001000110 : data_out = 24'b000000000000000100001000;
    16'b1111001001000111 : data_out = 24'b000000000000000100001001;
    16'b1111001001001000 : data_out = 24'b000000000000000100001001;
    16'b1111001001001001 : data_out = 24'b000000000000000100001001;
    16'b1111001001001010 : data_out = 24'b000000000000000100001001;
    16'b1111001001001011 : data_out = 24'b000000000000000100001010;
    16'b1111001001001100 : data_out = 24'b000000000000000100001010;
    16'b1111001001001101 : data_out = 24'b000000000000000100001010;
    16'b1111001001001110 : data_out = 24'b000000000000000100001010;
    16'b1111001001001111 : data_out = 24'b000000000000000100001011;
    16'b1111001001010000 : data_out = 24'b000000000000000100001011;
    16'b1111001001010001 : data_out = 24'b000000000000000100001011;
    16'b1111001001010010 : data_out = 24'b000000000000000100001100;
    16'b1111001001010011 : data_out = 24'b000000000000000100001100;
    16'b1111001001010100 : data_out = 24'b000000000000000100001100;
    16'b1111001001010101 : data_out = 24'b000000000000000100001100;
    16'b1111001001010110 : data_out = 24'b000000000000000100001101;
    16'b1111001001010111 : data_out = 24'b000000000000000100001101;
    16'b1111001001011000 : data_out = 24'b000000000000000100001101;
    16'b1111001001011001 : data_out = 24'b000000000000000100001101;
    16'b1111001001011010 : data_out = 24'b000000000000000100001110;
    16'b1111001001011011 : data_out = 24'b000000000000000100001110;
    16'b1111001001011100 : data_out = 24'b000000000000000100001110;
    16'b1111001001011101 : data_out = 24'b000000000000000100001110;
    16'b1111001001011110 : data_out = 24'b000000000000000100001111;
    16'b1111001001011111 : data_out = 24'b000000000000000100001111;
    16'b1111001001100000 : data_out = 24'b000000000000000100001111;
    16'b1111001001100001 : data_out = 24'b000000000000000100001111;
    16'b1111001001100010 : data_out = 24'b000000000000000100010000;
    16'b1111001001100011 : data_out = 24'b000000000000000100010000;
    16'b1111001001100100 : data_out = 24'b000000000000000100010000;
    16'b1111001001100101 : data_out = 24'b000000000000000100010001;
    16'b1111001001100110 : data_out = 24'b000000000000000100010001;
    16'b1111001001100111 : data_out = 24'b000000000000000100010001;
    16'b1111001001101000 : data_out = 24'b000000000000000100010001;
    16'b1111001001101001 : data_out = 24'b000000000000000100010010;
    16'b1111001001101010 : data_out = 24'b000000000000000100010010;
    16'b1111001001101011 : data_out = 24'b000000000000000100010010;
    16'b1111001001101100 : data_out = 24'b000000000000000100010010;
    16'b1111001001101101 : data_out = 24'b000000000000000100010011;
    16'b1111001001101110 : data_out = 24'b000000000000000100010011;
    16'b1111001001101111 : data_out = 24'b000000000000000100010011;
    16'b1111001001110000 : data_out = 24'b000000000000000100010011;
    16'b1111001001110001 : data_out = 24'b000000000000000100010100;
    16'b1111001001110010 : data_out = 24'b000000000000000100010100;
    16'b1111001001110011 : data_out = 24'b000000000000000100010100;
    16'b1111001001110100 : data_out = 24'b000000000000000100010101;
    16'b1111001001110101 : data_out = 24'b000000000000000100010101;
    16'b1111001001110110 : data_out = 24'b000000000000000100010101;
    16'b1111001001110111 : data_out = 24'b000000000000000100010101;
    16'b1111001001111000 : data_out = 24'b000000000000000100010110;
    16'b1111001001111001 : data_out = 24'b000000000000000100010110;
    16'b1111001001111010 : data_out = 24'b000000000000000100010110;
    16'b1111001001111011 : data_out = 24'b000000000000000100010110;
    16'b1111001001111100 : data_out = 24'b000000000000000100010111;
    16'b1111001001111101 : data_out = 24'b000000000000000100010111;
    16'b1111001001111110 : data_out = 24'b000000000000000100010111;
    16'b1111001001111111 : data_out = 24'b000000000000000100011000;
    16'b1111001010000000 : data_out = 24'b000000000000000100011000;
    16'b1111001010000001 : data_out = 24'b000000000000000100011000;
    16'b1111001010000010 : data_out = 24'b000000000000000100011000;
    16'b1111001010000011 : data_out = 24'b000000000000000100011001;
    16'b1111001010000100 : data_out = 24'b000000000000000100011001;
    16'b1111001010000101 : data_out = 24'b000000000000000100011001;
    16'b1111001010000110 : data_out = 24'b000000000000000100011001;
    16'b1111001010000111 : data_out = 24'b000000000000000100011010;
    16'b1111001010001000 : data_out = 24'b000000000000000100011010;
    16'b1111001010001001 : data_out = 24'b000000000000000100011010;
    16'b1111001010001010 : data_out = 24'b000000000000000100011011;
    16'b1111001010001011 : data_out = 24'b000000000000000100011011;
    16'b1111001010001100 : data_out = 24'b000000000000000100011011;
    16'b1111001010001101 : data_out = 24'b000000000000000100011011;
    16'b1111001010001110 : data_out = 24'b000000000000000100011100;
    16'b1111001010001111 : data_out = 24'b000000000000000100011100;
    16'b1111001010010000 : data_out = 24'b000000000000000100011100;
    16'b1111001010010001 : data_out = 24'b000000000000000100011101;
    16'b1111001010010010 : data_out = 24'b000000000000000100011101;
    16'b1111001010010011 : data_out = 24'b000000000000000100011101;
    16'b1111001010010100 : data_out = 24'b000000000000000100011101;
    16'b1111001010010101 : data_out = 24'b000000000000000100011110;
    16'b1111001010010110 : data_out = 24'b000000000000000100011110;
    16'b1111001010010111 : data_out = 24'b000000000000000100011110;
    16'b1111001010011000 : data_out = 24'b000000000000000100011110;
    16'b1111001010011001 : data_out = 24'b000000000000000100011111;
    16'b1111001010011010 : data_out = 24'b000000000000000100011111;
    16'b1111001010011011 : data_out = 24'b000000000000000100011111;
    16'b1111001010011100 : data_out = 24'b000000000000000100100000;
    16'b1111001010011101 : data_out = 24'b000000000000000100100000;
    16'b1111001010011110 : data_out = 24'b000000000000000100100000;
    16'b1111001010011111 : data_out = 24'b000000000000000100100000;
    16'b1111001010100000 : data_out = 24'b000000000000000100100001;
    16'b1111001010100001 : data_out = 24'b000000000000000100100001;
    16'b1111001010100010 : data_out = 24'b000000000000000100100001;
    16'b1111001010100011 : data_out = 24'b000000000000000100100010;
    16'b1111001010100100 : data_out = 24'b000000000000000100100010;
    16'b1111001010100101 : data_out = 24'b000000000000000100100010;
    16'b1111001010100110 : data_out = 24'b000000000000000100100010;
    16'b1111001010100111 : data_out = 24'b000000000000000100100011;
    16'b1111001010101000 : data_out = 24'b000000000000000100100011;
    16'b1111001010101001 : data_out = 24'b000000000000000100100011;
    16'b1111001010101010 : data_out = 24'b000000000000000100100100;
    16'b1111001010101011 : data_out = 24'b000000000000000100100100;
    16'b1111001010101100 : data_out = 24'b000000000000000100100100;
    16'b1111001010101101 : data_out = 24'b000000000000000100100100;
    16'b1111001010101110 : data_out = 24'b000000000000000100100101;
    16'b1111001010101111 : data_out = 24'b000000000000000100100101;
    16'b1111001010110000 : data_out = 24'b000000000000000100100101;
    16'b1111001010110001 : data_out = 24'b000000000000000100100110;
    16'b1111001010110010 : data_out = 24'b000000000000000100100110;
    16'b1111001010110011 : data_out = 24'b000000000000000100100110;
    16'b1111001010110100 : data_out = 24'b000000000000000100100110;
    16'b1111001010110101 : data_out = 24'b000000000000000100100111;
    16'b1111001010110110 : data_out = 24'b000000000000000100100111;
    16'b1111001010110111 : data_out = 24'b000000000000000100100111;
    16'b1111001010111000 : data_out = 24'b000000000000000100101000;
    16'b1111001010111001 : data_out = 24'b000000000000000100101000;
    16'b1111001010111010 : data_out = 24'b000000000000000100101000;
    16'b1111001010111011 : data_out = 24'b000000000000000100101000;
    16'b1111001010111100 : data_out = 24'b000000000000000100101001;
    16'b1111001010111101 : data_out = 24'b000000000000000100101001;
    16'b1111001010111110 : data_out = 24'b000000000000000100101001;
    16'b1111001010111111 : data_out = 24'b000000000000000100101010;
    16'b1111001011000000 : data_out = 24'b000000000000000100101010;
    16'b1111001011000001 : data_out = 24'b000000000000000100101010;
    16'b1111001011000010 : data_out = 24'b000000000000000100101010;
    16'b1111001011000011 : data_out = 24'b000000000000000100101011;
    16'b1111001011000100 : data_out = 24'b000000000000000100101011;
    16'b1111001011000101 : data_out = 24'b000000000000000100101011;
    16'b1111001011000110 : data_out = 24'b000000000000000100101100;
    16'b1111001011000111 : data_out = 24'b000000000000000100101100;
    16'b1111001011001000 : data_out = 24'b000000000000000100101100;
    16'b1111001011001001 : data_out = 24'b000000000000000100101101;
    16'b1111001011001010 : data_out = 24'b000000000000000100101101;
    16'b1111001011001011 : data_out = 24'b000000000000000100101101;
    16'b1111001011001100 : data_out = 24'b000000000000000100101101;
    16'b1111001011001101 : data_out = 24'b000000000000000100101110;
    16'b1111001011001110 : data_out = 24'b000000000000000100101110;
    16'b1111001011001111 : data_out = 24'b000000000000000100101110;
    16'b1111001011010000 : data_out = 24'b000000000000000100101111;
    16'b1111001011010001 : data_out = 24'b000000000000000100101111;
    16'b1111001011010010 : data_out = 24'b000000000000000100101111;
    16'b1111001011010011 : data_out = 24'b000000000000000100101111;
    16'b1111001011010100 : data_out = 24'b000000000000000100110000;
    16'b1111001011010101 : data_out = 24'b000000000000000100110000;
    16'b1111001011010110 : data_out = 24'b000000000000000100110000;
    16'b1111001011010111 : data_out = 24'b000000000000000100110001;
    16'b1111001011011000 : data_out = 24'b000000000000000100110001;
    16'b1111001011011001 : data_out = 24'b000000000000000100110001;
    16'b1111001011011010 : data_out = 24'b000000000000000100110010;
    16'b1111001011011011 : data_out = 24'b000000000000000100110010;
    16'b1111001011011100 : data_out = 24'b000000000000000100110010;
    16'b1111001011011101 : data_out = 24'b000000000000000100110010;
    16'b1111001011011110 : data_out = 24'b000000000000000100110011;
    16'b1111001011011111 : data_out = 24'b000000000000000100110011;
    16'b1111001011100000 : data_out = 24'b000000000000000100110011;
    16'b1111001011100001 : data_out = 24'b000000000000000100110100;
    16'b1111001011100010 : data_out = 24'b000000000000000100110100;
    16'b1111001011100011 : data_out = 24'b000000000000000100110100;
    16'b1111001011100100 : data_out = 24'b000000000000000100110101;
    16'b1111001011100101 : data_out = 24'b000000000000000100110101;
    16'b1111001011100110 : data_out = 24'b000000000000000100110101;
    16'b1111001011100111 : data_out = 24'b000000000000000100110101;
    16'b1111001011101000 : data_out = 24'b000000000000000100110110;
    16'b1111001011101001 : data_out = 24'b000000000000000100110110;
    16'b1111001011101010 : data_out = 24'b000000000000000100110110;
    16'b1111001011101011 : data_out = 24'b000000000000000100110111;
    16'b1111001011101100 : data_out = 24'b000000000000000100110111;
    16'b1111001011101101 : data_out = 24'b000000000000000100110111;
    16'b1111001011101110 : data_out = 24'b000000000000000100111000;
    16'b1111001011101111 : data_out = 24'b000000000000000100111000;
    16'b1111001011110000 : data_out = 24'b000000000000000100111000;
    16'b1111001011110001 : data_out = 24'b000000000000000100111001;
    16'b1111001011110010 : data_out = 24'b000000000000000100111001;
    16'b1111001011110011 : data_out = 24'b000000000000000100111001;
    16'b1111001011110100 : data_out = 24'b000000000000000100111001;
    16'b1111001011110101 : data_out = 24'b000000000000000100111010;
    16'b1111001011110110 : data_out = 24'b000000000000000100111010;
    16'b1111001011110111 : data_out = 24'b000000000000000100111010;
    16'b1111001011111000 : data_out = 24'b000000000000000100111011;
    16'b1111001011111001 : data_out = 24'b000000000000000100111011;
    16'b1111001011111010 : data_out = 24'b000000000000000100111011;
    16'b1111001011111011 : data_out = 24'b000000000000000100111100;
    16'b1111001011111100 : data_out = 24'b000000000000000100111100;
    16'b1111001011111101 : data_out = 24'b000000000000000100111100;
    16'b1111001011111110 : data_out = 24'b000000000000000100111101;
    16'b1111001011111111 : data_out = 24'b000000000000000100111101;
    16'b1111001100000000 : data_out = 24'b000000000000000100111101;
    16'b1111001100000001 : data_out = 24'b000000000000000100111101;
    16'b1111001100000010 : data_out = 24'b000000000000000100111110;
    16'b1111001100000011 : data_out = 24'b000000000000000100111110;
    16'b1111001100000100 : data_out = 24'b000000000000000100111110;
    16'b1111001100000101 : data_out = 24'b000000000000000100111111;
    16'b1111001100000110 : data_out = 24'b000000000000000100111111;
    16'b1111001100000111 : data_out = 24'b000000000000000100111111;
    16'b1111001100001000 : data_out = 24'b000000000000000101000000;
    16'b1111001100001001 : data_out = 24'b000000000000000101000000;
    16'b1111001100001010 : data_out = 24'b000000000000000101000000;
    16'b1111001100001011 : data_out = 24'b000000000000000101000001;
    16'b1111001100001100 : data_out = 24'b000000000000000101000001;
    16'b1111001100001101 : data_out = 24'b000000000000000101000001;
    16'b1111001100001110 : data_out = 24'b000000000000000101000010;
    16'b1111001100001111 : data_out = 24'b000000000000000101000010;
    16'b1111001100010000 : data_out = 24'b000000000000000101000010;
    16'b1111001100010001 : data_out = 24'b000000000000000101000010;
    16'b1111001100010010 : data_out = 24'b000000000000000101000011;
    16'b1111001100010011 : data_out = 24'b000000000000000101000011;
    16'b1111001100010100 : data_out = 24'b000000000000000101000011;
    16'b1111001100010101 : data_out = 24'b000000000000000101000100;
    16'b1111001100010110 : data_out = 24'b000000000000000101000100;
    16'b1111001100010111 : data_out = 24'b000000000000000101000100;
    16'b1111001100011000 : data_out = 24'b000000000000000101000101;
    16'b1111001100011001 : data_out = 24'b000000000000000101000101;
    16'b1111001100011010 : data_out = 24'b000000000000000101000101;
    16'b1111001100011011 : data_out = 24'b000000000000000101000110;
    16'b1111001100011100 : data_out = 24'b000000000000000101000110;
    16'b1111001100011101 : data_out = 24'b000000000000000101000110;
    16'b1111001100011110 : data_out = 24'b000000000000000101000111;
    16'b1111001100011111 : data_out = 24'b000000000000000101000111;
    16'b1111001100100000 : data_out = 24'b000000000000000101000111;
    16'b1111001100100001 : data_out = 24'b000000000000000101001000;
    16'b1111001100100010 : data_out = 24'b000000000000000101001000;
    16'b1111001100100011 : data_out = 24'b000000000000000101001000;
    16'b1111001100100100 : data_out = 24'b000000000000000101001001;
    16'b1111001100100101 : data_out = 24'b000000000000000101001001;
    16'b1111001100100110 : data_out = 24'b000000000000000101001001;
    16'b1111001100100111 : data_out = 24'b000000000000000101001001;
    16'b1111001100101000 : data_out = 24'b000000000000000101001010;
    16'b1111001100101001 : data_out = 24'b000000000000000101001010;
    16'b1111001100101010 : data_out = 24'b000000000000000101001010;
    16'b1111001100101011 : data_out = 24'b000000000000000101001011;
    16'b1111001100101100 : data_out = 24'b000000000000000101001011;
    16'b1111001100101101 : data_out = 24'b000000000000000101001011;
    16'b1111001100101110 : data_out = 24'b000000000000000101001100;
    16'b1111001100101111 : data_out = 24'b000000000000000101001100;
    16'b1111001100110000 : data_out = 24'b000000000000000101001100;
    16'b1111001100110001 : data_out = 24'b000000000000000101001101;
    16'b1111001100110010 : data_out = 24'b000000000000000101001101;
    16'b1111001100110011 : data_out = 24'b000000000000000101001101;
    16'b1111001100110100 : data_out = 24'b000000000000000101001110;
    16'b1111001100110101 : data_out = 24'b000000000000000101001110;
    16'b1111001100110110 : data_out = 24'b000000000000000101001110;
    16'b1111001100110111 : data_out = 24'b000000000000000101001111;
    16'b1111001100111000 : data_out = 24'b000000000000000101001111;
    16'b1111001100111001 : data_out = 24'b000000000000000101001111;
    16'b1111001100111010 : data_out = 24'b000000000000000101010000;
    16'b1111001100111011 : data_out = 24'b000000000000000101010000;
    16'b1111001100111100 : data_out = 24'b000000000000000101010000;
    16'b1111001100111101 : data_out = 24'b000000000000000101010001;
    16'b1111001100111110 : data_out = 24'b000000000000000101010001;
    16'b1111001100111111 : data_out = 24'b000000000000000101010001;
    16'b1111001101000000 : data_out = 24'b000000000000000101010010;
    16'b1111001101000001 : data_out = 24'b000000000000000101010010;
    16'b1111001101000010 : data_out = 24'b000000000000000101010010;
    16'b1111001101000011 : data_out = 24'b000000000000000101010011;
    16'b1111001101000100 : data_out = 24'b000000000000000101010011;
    16'b1111001101000101 : data_out = 24'b000000000000000101010011;
    16'b1111001101000110 : data_out = 24'b000000000000000101010100;
    16'b1111001101000111 : data_out = 24'b000000000000000101010100;
    16'b1111001101001000 : data_out = 24'b000000000000000101010100;
    16'b1111001101001001 : data_out = 24'b000000000000000101010101;
    16'b1111001101001010 : data_out = 24'b000000000000000101010101;
    16'b1111001101001011 : data_out = 24'b000000000000000101010101;
    16'b1111001101001100 : data_out = 24'b000000000000000101010110;
    16'b1111001101001101 : data_out = 24'b000000000000000101010110;
    16'b1111001101001110 : data_out = 24'b000000000000000101010110;
    16'b1111001101001111 : data_out = 24'b000000000000000101010111;
    16'b1111001101010000 : data_out = 24'b000000000000000101010111;
    16'b1111001101010001 : data_out = 24'b000000000000000101010111;
    16'b1111001101010010 : data_out = 24'b000000000000000101011000;
    16'b1111001101010011 : data_out = 24'b000000000000000101011000;
    16'b1111001101010100 : data_out = 24'b000000000000000101011000;
    16'b1111001101010101 : data_out = 24'b000000000000000101011001;
    16'b1111001101010110 : data_out = 24'b000000000000000101011001;
    16'b1111001101010111 : data_out = 24'b000000000000000101011001;
    16'b1111001101011000 : data_out = 24'b000000000000000101011010;
    16'b1111001101011001 : data_out = 24'b000000000000000101011010;
    16'b1111001101011010 : data_out = 24'b000000000000000101011010;
    16'b1111001101011011 : data_out = 24'b000000000000000101011011;
    16'b1111001101011100 : data_out = 24'b000000000000000101011011;
    16'b1111001101011101 : data_out = 24'b000000000000000101011011;
    16'b1111001101011110 : data_out = 24'b000000000000000101011100;
    16'b1111001101011111 : data_out = 24'b000000000000000101011100;
    16'b1111001101100000 : data_out = 24'b000000000000000101011100;
    16'b1111001101100001 : data_out = 24'b000000000000000101011101;
    16'b1111001101100010 : data_out = 24'b000000000000000101011101;
    16'b1111001101100011 : data_out = 24'b000000000000000101011101;
    16'b1111001101100100 : data_out = 24'b000000000000000101011110;
    16'b1111001101100101 : data_out = 24'b000000000000000101011110;
    16'b1111001101100110 : data_out = 24'b000000000000000101011110;
    16'b1111001101100111 : data_out = 24'b000000000000000101011111;
    16'b1111001101101000 : data_out = 24'b000000000000000101011111;
    16'b1111001101101001 : data_out = 24'b000000000000000101011111;
    16'b1111001101101010 : data_out = 24'b000000000000000101100000;
    16'b1111001101101011 : data_out = 24'b000000000000000101100000;
    16'b1111001101101100 : data_out = 24'b000000000000000101100000;
    16'b1111001101101101 : data_out = 24'b000000000000000101100001;
    16'b1111001101101110 : data_out = 24'b000000000000000101100001;
    16'b1111001101101111 : data_out = 24'b000000000000000101100010;
    16'b1111001101110000 : data_out = 24'b000000000000000101100010;
    16'b1111001101110001 : data_out = 24'b000000000000000101100010;
    16'b1111001101110010 : data_out = 24'b000000000000000101100011;
    16'b1111001101110011 : data_out = 24'b000000000000000101100011;
    16'b1111001101110100 : data_out = 24'b000000000000000101100011;
    16'b1111001101110101 : data_out = 24'b000000000000000101100100;
    16'b1111001101110110 : data_out = 24'b000000000000000101100100;
    16'b1111001101110111 : data_out = 24'b000000000000000101100100;
    16'b1111001101111000 : data_out = 24'b000000000000000101100101;
    16'b1111001101111001 : data_out = 24'b000000000000000101100101;
    16'b1111001101111010 : data_out = 24'b000000000000000101100101;
    16'b1111001101111011 : data_out = 24'b000000000000000101100110;
    16'b1111001101111100 : data_out = 24'b000000000000000101100110;
    16'b1111001101111101 : data_out = 24'b000000000000000101100110;
    16'b1111001101111110 : data_out = 24'b000000000000000101100111;
    16'b1111001101111111 : data_out = 24'b000000000000000101100111;
    16'b1111001110000000 : data_out = 24'b000000000000000101100111;
    16'b1111001110000001 : data_out = 24'b000000000000000101101000;
    16'b1111001110000010 : data_out = 24'b000000000000000101101000;
    16'b1111001110000011 : data_out = 24'b000000000000000101101000;
    16'b1111001110000100 : data_out = 24'b000000000000000101101001;
    16'b1111001110000101 : data_out = 24'b000000000000000101101001;
    16'b1111001110000110 : data_out = 24'b000000000000000101101010;
    16'b1111001110000111 : data_out = 24'b000000000000000101101010;
    16'b1111001110001000 : data_out = 24'b000000000000000101101010;
    16'b1111001110001001 : data_out = 24'b000000000000000101101011;
    16'b1111001110001010 : data_out = 24'b000000000000000101101011;
    16'b1111001110001011 : data_out = 24'b000000000000000101101011;
    16'b1111001110001100 : data_out = 24'b000000000000000101101100;
    16'b1111001110001101 : data_out = 24'b000000000000000101101100;
    16'b1111001110001110 : data_out = 24'b000000000000000101101100;
    16'b1111001110001111 : data_out = 24'b000000000000000101101101;
    16'b1111001110010000 : data_out = 24'b000000000000000101101101;
    16'b1111001110010001 : data_out = 24'b000000000000000101101101;
    16'b1111001110010010 : data_out = 24'b000000000000000101101110;
    16'b1111001110010011 : data_out = 24'b000000000000000101101110;
    16'b1111001110010100 : data_out = 24'b000000000000000101101111;
    16'b1111001110010101 : data_out = 24'b000000000000000101101111;
    16'b1111001110010110 : data_out = 24'b000000000000000101101111;
    16'b1111001110010111 : data_out = 24'b000000000000000101110000;
    16'b1111001110011000 : data_out = 24'b000000000000000101110000;
    16'b1111001110011001 : data_out = 24'b000000000000000101110000;
    16'b1111001110011010 : data_out = 24'b000000000000000101110001;
    16'b1111001110011011 : data_out = 24'b000000000000000101110001;
    16'b1111001110011100 : data_out = 24'b000000000000000101110001;
    16'b1111001110011101 : data_out = 24'b000000000000000101110010;
    16'b1111001110011110 : data_out = 24'b000000000000000101110010;
    16'b1111001110011111 : data_out = 24'b000000000000000101110010;
    16'b1111001110100000 : data_out = 24'b000000000000000101110011;
    16'b1111001110100001 : data_out = 24'b000000000000000101110011;
    16'b1111001110100010 : data_out = 24'b000000000000000101110100;
    16'b1111001110100011 : data_out = 24'b000000000000000101110100;
    16'b1111001110100100 : data_out = 24'b000000000000000101110100;
    16'b1111001110100101 : data_out = 24'b000000000000000101110101;
    16'b1111001110100110 : data_out = 24'b000000000000000101110101;
    16'b1111001110100111 : data_out = 24'b000000000000000101110101;
    16'b1111001110101000 : data_out = 24'b000000000000000101110110;
    16'b1111001110101001 : data_out = 24'b000000000000000101110110;
    16'b1111001110101010 : data_out = 24'b000000000000000101110111;
    16'b1111001110101011 : data_out = 24'b000000000000000101110111;
    16'b1111001110101100 : data_out = 24'b000000000000000101110111;
    16'b1111001110101101 : data_out = 24'b000000000000000101111000;
    16'b1111001110101110 : data_out = 24'b000000000000000101111000;
    16'b1111001110101111 : data_out = 24'b000000000000000101111000;
    16'b1111001110110000 : data_out = 24'b000000000000000101111001;
    16'b1111001110110001 : data_out = 24'b000000000000000101111001;
    16'b1111001110110010 : data_out = 24'b000000000000000101111001;
    16'b1111001110110011 : data_out = 24'b000000000000000101111010;
    16'b1111001110110100 : data_out = 24'b000000000000000101111010;
    16'b1111001110110101 : data_out = 24'b000000000000000101111011;
    16'b1111001110110110 : data_out = 24'b000000000000000101111011;
    16'b1111001110110111 : data_out = 24'b000000000000000101111011;
    16'b1111001110111000 : data_out = 24'b000000000000000101111100;
    16'b1111001110111001 : data_out = 24'b000000000000000101111100;
    16'b1111001110111010 : data_out = 24'b000000000000000101111100;
    16'b1111001110111011 : data_out = 24'b000000000000000101111101;
    16'b1111001110111100 : data_out = 24'b000000000000000101111101;
    16'b1111001110111101 : data_out = 24'b000000000000000101111110;
    16'b1111001110111110 : data_out = 24'b000000000000000101111110;
    16'b1111001110111111 : data_out = 24'b000000000000000101111110;
    16'b1111001111000000 : data_out = 24'b000000000000000101111111;
    16'b1111001111000001 : data_out = 24'b000000000000000101111111;
    16'b1111001111000010 : data_out = 24'b000000000000000101111111;
    16'b1111001111000011 : data_out = 24'b000000000000000110000000;
    16'b1111001111000100 : data_out = 24'b000000000000000110000000;
    16'b1111001111000101 : data_out = 24'b000000000000000110000001;
    16'b1111001111000110 : data_out = 24'b000000000000000110000001;
    16'b1111001111000111 : data_out = 24'b000000000000000110000001;
    16'b1111001111001000 : data_out = 24'b000000000000000110000010;
    16'b1111001111001001 : data_out = 24'b000000000000000110000010;
    16'b1111001111001010 : data_out = 24'b000000000000000110000010;
    16'b1111001111001011 : data_out = 24'b000000000000000110000011;
    16'b1111001111001100 : data_out = 24'b000000000000000110000011;
    16'b1111001111001101 : data_out = 24'b000000000000000110000100;
    16'b1111001111001110 : data_out = 24'b000000000000000110000100;
    16'b1111001111001111 : data_out = 24'b000000000000000110000100;
    16'b1111001111010000 : data_out = 24'b000000000000000110000101;
    16'b1111001111010001 : data_out = 24'b000000000000000110000101;
    16'b1111001111010010 : data_out = 24'b000000000000000110000101;
    16'b1111001111010011 : data_out = 24'b000000000000000110000110;
    16'b1111001111010100 : data_out = 24'b000000000000000110000110;
    16'b1111001111010101 : data_out = 24'b000000000000000110000111;
    16'b1111001111010110 : data_out = 24'b000000000000000110000111;
    16'b1111001111010111 : data_out = 24'b000000000000000110000111;
    16'b1111001111011000 : data_out = 24'b000000000000000110001000;
    16'b1111001111011001 : data_out = 24'b000000000000000110001000;
    16'b1111001111011010 : data_out = 24'b000000000000000110001000;
    16'b1111001111011011 : data_out = 24'b000000000000000110001001;
    16'b1111001111011100 : data_out = 24'b000000000000000110001001;
    16'b1111001111011101 : data_out = 24'b000000000000000110001010;
    16'b1111001111011110 : data_out = 24'b000000000000000110001010;
    16'b1111001111011111 : data_out = 24'b000000000000000110001010;
    16'b1111001111100000 : data_out = 24'b000000000000000110001011;
    16'b1111001111100001 : data_out = 24'b000000000000000110001011;
    16'b1111001111100010 : data_out = 24'b000000000000000110001100;
    16'b1111001111100011 : data_out = 24'b000000000000000110001100;
    16'b1111001111100100 : data_out = 24'b000000000000000110001100;
    16'b1111001111100101 : data_out = 24'b000000000000000110001101;
    16'b1111001111100110 : data_out = 24'b000000000000000110001101;
    16'b1111001111100111 : data_out = 24'b000000000000000110001110;
    16'b1111001111101000 : data_out = 24'b000000000000000110001110;
    16'b1111001111101001 : data_out = 24'b000000000000000110001110;
    16'b1111001111101010 : data_out = 24'b000000000000000110001111;
    16'b1111001111101011 : data_out = 24'b000000000000000110001111;
    16'b1111001111101100 : data_out = 24'b000000000000000110001111;
    16'b1111001111101101 : data_out = 24'b000000000000000110010000;
    16'b1111001111101110 : data_out = 24'b000000000000000110010000;
    16'b1111001111101111 : data_out = 24'b000000000000000110010001;
    16'b1111001111110000 : data_out = 24'b000000000000000110010001;
    16'b1111001111110001 : data_out = 24'b000000000000000110010001;
    16'b1111001111110010 : data_out = 24'b000000000000000110010010;
    16'b1111001111110011 : data_out = 24'b000000000000000110010010;
    16'b1111001111110100 : data_out = 24'b000000000000000110010011;
    16'b1111001111110101 : data_out = 24'b000000000000000110010011;
    16'b1111001111110110 : data_out = 24'b000000000000000110010011;
    16'b1111001111110111 : data_out = 24'b000000000000000110010100;
    16'b1111001111111000 : data_out = 24'b000000000000000110010100;
    16'b1111001111111001 : data_out = 24'b000000000000000110010101;
    16'b1111001111111010 : data_out = 24'b000000000000000110010101;
    16'b1111001111111011 : data_out = 24'b000000000000000110010101;
    16'b1111001111111100 : data_out = 24'b000000000000000110010110;
    16'b1111001111111101 : data_out = 24'b000000000000000110010110;
    16'b1111001111111110 : data_out = 24'b000000000000000110010111;
    16'b1111001111111111 : data_out = 24'b000000000000000110010111;
    16'b1111010000000000 : data_out = 24'b000000000000000110010111;
    16'b1111010000000001 : data_out = 24'b000000000000000110011000;
    16'b1111010000000010 : data_out = 24'b000000000000000110011000;
    16'b1111010000000011 : data_out = 24'b000000000000000110011001;
    16'b1111010000000100 : data_out = 24'b000000000000000110011001;
    16'b1111010000000101 : data_out = 24'b000000000000000110011001;
    16'b1111010000000110 : data_out = 24'b000000000000000110011010;
    16'b1111010000000111 : data_out = 24'b000000000000000110011010;
    16'b1111010000001000 : data_out = 24'b000000000000000110011011;
    16'b1111010000001001 : data_out = 24'b000000000000000110011011;
    16'b1111010000001010 : data_out = 24'b000000000000000110011011;
    16'b1111010000001011 : data_out = 24'b000000000000000110011100;
    16'b1111010000001100 : data_out = 24'b000000000000000110011100;
    16'b1111010000001101 : data_out = 24'b000000000000000110011101;
    16'b1111010000001110 : data_out = 24'b000000000000000110011101;
    16'b1111010000001111 : data_out = 24'b000000000000000110011101;
    16'b1111010000010000 : data_out = 24'b000000000000000110011110;
    16'b1111010000010001 : data_out = 24'b000000000000000110011110;
    16'b1111010000010010 : data_out = 24'b000000000000000110011111;
    16'b1111010000010011 : data_out = 24'b000000000000000110011111;
    16'b1111010000010100 : data_out = 24'b000000000000000110011111;
    16'b1111010000010101 : data_out = 24'b000000000000000110100000;
    16'b1111010000010110 : data_out = 24'b000000000000000110100000;
    16'b1111010000010111 : data_out = 24'b000000000000000110100001;
    16'b1111010000011000 : data_out = 24'b000000000000000110100001;
    16'b1111010000011001 : data_out = 24'b000000000000000110100001;
    16'b1111010000011010 : data_out = 24'b000000000000000110100010;
    16'b1111010000011011 : data_out = 24'b000000000000000110100010;
    16'b1111010000011100 : data_out = 24'b000000000000000110100011;
    16'b1111010000011101 : data_out = 24'b000000000000000110100011;
    16'b1111010000011110 : data_out = 24'b000000000000000110100011;
    16'b1111010000011111 : data_out = 24'b000000000000000110100100;
    16'b1111010000100000 : data_out = 24'b000000000000000110100100;
    16'b1111010000100001 : data_out = 24'b000000000000000110100101;
    16'b1111010000100010 : data_out = 24'b000000000000000110100101;
    16'b1111010000100011 : data_out = 24'b000000000000000110100110;
    16'b1111010000100100 : data_out = 24'b000000000000000110100110;
    16'b1111010000100101 : data_out = 24'b000000000000000110100110;
    16'b1111010000100110 : data_out = 24'b000000000000000110100111;
    16'b1111010000100111 : data_out = 24'b000000000000000110100111;
    16'b1111010000101000 : data_out = 24'b000000000000000110101000;
    16'b1111010000101001 : data_out = 24'b000000000000000110101000;
    16'b1111010000101010 : data_out = 24'b000000000000000110101000;
    16'b1111010000101011 : data_out = 24'b000000000000000110101001;
    16'b1111010000101100 : data_out = 24'b000000000000000110101001;
    16'b1111010000101101 : data_out = 24'b000000000000000110101010;
    16'b1111010000101110 : data_out = 24'b000000000000000110101010;
    16'b1111010000101111 : data_out = 24'b000000000000000110101011;
    16'b1111010000110000 : data_out = 24'b000000000000000110101011;
    16'b1111010000110001 : data_out = 24'b000000000000000110101011;
    16'b1111010000110010 : data_out = 24'b000000000000000110101100;
    16'b1111010000110011 : data_out = 24'b000000000000000110101100;
    16'b1111010000110100 : data_out = 24'b000000000000000110101101;
    16'b1111010000110101 : data_out = 24'b000000000000000110101101;
    16'b1111010000110110 : data_out = 24'b000000000000000110101101;
    16'b1111010000110111 : data_out = 24'b000000000000000110101110;
    16'b1111010000111000 : data_out = 24'b000000000000000110101110;
    16'b1111010000111001 : data_out = 24'b000000000000000110101111;
    16'b1111010000111010 : data_out = 24'b000000000000000110101111;
    16'b1111010000111011 : data_out = 24'b000000000000000110110000;
    16'b1111010000111100 : data_out = 24'b000000000000000110110000;
    16'b1111010000111101 : data_out = 24'b000000000000000110110000;
    16'b1111010000111110 : data_out = 24'b000000000000000110110001;
    16'b1111010000111111 : data_out = 24'b000000000000000110110001;
    16'b1111010001000000 : data_out = 24'b000000000000000110110010;
    16'b1111010001000001 : data_out = 24'b000000000000000110110010;
    16'b1111010001000010 : data_out = 24'b000000000000000110110011;
    16'b1111010001000011 : data_out = 24'b000000000000000110110011;
    16'b1111010001000100 : data_out = 24'b000000000000000110110011;
    16'b1111010001000101 : data_out = 24'b000000000000000110110100;
    16'b1111010001000110 : data_out = 24'b000000000000000110110100;
    16'b1111010001000111 : data_out = 24'b000000000000000110110101;
    16'b1111010001001000 : data_out = 24'b000000000000000110110101;
    16'b1111010001001001 : data_out = 24'b000000000000000110110101;
    16'b1111010001001010 : data_out = 24'b000000000000000110110110;
    16'b1111010001001011 : data_out = 24'b000000000000000110110110;
    16'b1111010001001100 : data_out = 24'b000000000000000110110111;
    16'b1111010001001101 : data_out = 24'b000000000000000110110111;
    16'b1111010001001110 : data_out = 24'b000000000000000110111000;
    16'b1111010001001111 : data_out = 24'b000000000000000110111000;
    16'b1111010001010000 : data_out = 24'b000000000000000110111000;
    16'b1111010001010001 : data_out = 24'b000000000000000110111001;
    16'b1111010001010010 : data_out = 24'b000000000000000110111001;
    16'b1111010001010011 : data_out = 24'b000000000000000110111010;
    16'b1111010001010100 : data_out = 24'b000000000000000110111010;
    16'b1111010001010101 : data_out = 24'b000000000000000110111011;
    16'b1111010001010110 : data_out = 24'b000000000000000110111011;
    16'b1111010001010111 : data_out = 24'b000000000000000110111100;
    16'b1111010001011000 : data_out = 24'b000000000000000110111100;
    16'b1111010001011001 : data_out = 24'b000000000000000110111100;
    16'b1111010001011010 : data_out = 24'b000000000000000110111101;
    16'b1111010001011011 : data_out = 24'b000000000000000110111101;
    16'b1111010001011100 : data_out = 24'b000000000000000110111110;
    16'b1111010001011101 : data_out = 24'b000000000000000110111110;
    16'b1111010001011110 : data_out = 24'b000000000000000110111111;
    16'b1111010001011111 : data_out = 24'b000000000000000110111111;
    16'b1111010001100000 : data_out = 24'b000000000000000110111111;
    16'b1111010001100001 : data_out = 24'b000000000000000111000000;
    16'b1111010001100010 : data_out = 24'b000000000000000111000000;
    16'b1111010001100011 : data_out = 24'b000000000000000111000001;
    16'b1111010001100100 : data_out = 24'b000000000000000111000001;
    16'b1111010001100101 : data_out = 24'b000000000000000111000010;
    16'b1111010001100110 : data_out = 24'b000000000000000111000010;
    16'b1111010001100111 : data_out = 24'b000000000000000111000011;
    16'b1111010001101000 : data_out = 24'b000000000000000111000011;
    16'b1111010001101001 : data_out = 24'b000000000000000111000011;
    16'b1111010001101010 : data_out = 24'b000000000000000111000100;
    16'b1111010001101011 : data_out = 24'b000000000000000111000100;
    16'b1111010001101100 : data_out = 24'b000000000000000111000101;
    16'b1111010001101101 : data_out = 24'b000000000000000111000101;
    16'b1111010001101110 : data_out = 24'b000000000000000111000110;
    16'b1111010001101111 : data_out = 24'b000000000000000111000110;
    16'b1111010001110000 : data_out = 24'b000000000000000111000110;
    16'b1111010001110001 : data_out = 24'b000000000000000111000111;
    16'b1111010001110010 : data_out = 24'b000000000000000111000111;
    16'b1111010001110011 : data_out = 24'b000000000000000111001000;
    16'b1111010001110100 : data_out = 24'b000000000000000111001000;
    16'b1111010001110101 : data_out = 24'b000000000000000111001001;
    16'b1111010001110110 : data_out = 24'b000000000000000111001001;
    16'b1111010001110111 : data_out = 24'b000000000000000111001010;
    16'b1111010001111000 : data_out = 24'b000000000000000111001010;
    16'b1111010001111001 : data_out = 24'b000000000000000111001011;
    16'b1111010001111010 : data_out = 24'b000000000000000111001011;
    16'b1111010001111011 : data_out = 24'b000000000000000111001011;
    16'b1111010001111100 : data_out = 24'b000000000000000111001100;
    16'b1111010001111101 : data_out = 24'b000000000000000111001100;
    16'b1111010001111110 : data_out = 24'b000000000000000111001101;
    16'b1111010001111111 : data_out = 24'b000000000000000111001101;
    16'b1111010010000000 : data_out = 24'b000000000000000111001110;
    16'b1111010010000001 : data_out = 24'b000000000000000111001110;
    16'b1111010010000010 : data_out = 24'b000000000000000111001111;
    16'b1111010010000011 : data_out = 24'b000000000000000111001111;
    16'b1111010010000100 : data_out = 24'b000000000000000111001111;
    16'b1111010010000101 : data_out = 24'b000000000000000111010000;
    16'b1111010010000110 : data_out = 24'b000000000000000111010000;
    16'b1111010010000111 : data_out = 24'b000000000000000111010001;
    16'b1111010010001000 : data_out = 24'b000000000000000111010001;
    16'b1111010010001001 : data_out = 24'b000000000000000111010010;
    16'b1111010010001010 : data_out = 24'b000000000000000111010010;
    16'b1111010010001011 : data_out = 24'b000000000000000111010011;
    16'b1111010010001100 : data_out = 24'b000000000000000111010011;
    16'b1111010010001101 : data_out = 24'b000000000000000111010100;
    16'b1111010010001110 : data_out = 24'b000000000000000111010100;
    16'b1111010010001111 : data_out = 24'b000000000000000111010100;
    16'b1111010010010000 : data_out = 24'b000000000000000111010101;
    16'b1111010010010001 : data_out = 24'b000000000000000111010101;
    16'b1111010010010010 : data_out = 24'b000000000000000111010110;
    16'b1111010010010011 : data_out = 24'b000000000000000111010110;
    16'b1111010010010100 : data_out = 24'b000000000000000111010111;
    16'b1111010010010101 : data_out = 24'b000000000000000111010111;
    16'b1111010010010110 : data_out = 24'b000000000000000111011000;
    16'b1111010010010111 : data_out = 24'b000000000000000111011000;
    16'b1111010010011000 : data_out = 24'b000000000000000111011001;
    16'b1111010010011001 : data_out = 24'b000000000000000111011001;
    16'b1111010010011010 : data_out = 24'b000000000000000111011010;
    16'b1111010010011011 : data_out = 24'b000000000000000111011010;
    16'b1111010010011100 : data_out = 24'b000000000000000111011010;
    16'b1111010010011101 : data_out = 24'b000000000000000111011011;
    16'b1111010010011110 : data_out = 24'b000000000000000111011011;
    16'b1111010010011111 : data_out = 24'b000000000000000111011100;
    16'b1111010010100000 : data_out = 24'b000000000000000111011100;
    16'b1111010010100001 : data_out = 24'b000000000000000111011101;
    16'b1111010010100010 : data_out = 24'b000000000000000111011101;
    16'b1111010010100011 : data_out = 24'b000000000000000111011110;
    16'b1111010010100100 : data_out = 24'b000000000000000111011110;
    16'b1111010010100101 : data_out = 24'b000000000000000111011111;
    16'b1111010010100110 : data_out = 24'b000000000000000111011111;
    16'b1111010010100111 : data_out = 24'b000000000000000111100000;
    16'b1111010010101000 : data_out = 24'b000000000000000111100000;
    16'b1111010010101001 : data_out = 24'b000000000000000111100001;
    16'b1111010010101010 : data_out = 24'b000000000000000111100001;
    16'b1111010010101011 : data_out = 24'b000000000000000111100001;
    16'b1111010010101100 : data_out = 24'b000000000000000111100010;
    16'b1111010010101101 : data_out = 24'b000000000000000111100010;
    16'b1111010010101110 : data_out = 24'b000000000000000111100011;
    16'b1111010010101111 : data_out = 24'b000000000000000111100011;
    16'b1111010010110000 : data_out = 24'b000000000000000111100100;
    16'b1111010010110001 : data_out = 24'b000000000000000111100100;
    16'b1111010010110010 : data_out = 24'b000000000000000111100101;
    16'b1111010010110011 : data_out = 24'b000000000000000111100101;
    16'b1111010010110100 : data_out = 24'b000000000000000111100110;
    16'b1111010010110101 : data_out = 24'b000000000000000111100110;
    16'b1111010010110110 : data_out = 24'b000000000000000111100111;
    16'b1111010010110111 : data_out = 24'b000000000000000111100111;
    16'b1111010010111000 : data_out = 24'b000000000000000111101000;
    16'b1111010010111001 : data_out = 24'b000000000000000111101000;
    16'b1111010010111010 : data_out = 24'b000000000000000111101001;
    16'b1111010010111011 : data_out = 24'b000000000000000111101001;
    16'b1111010010111100 : data_out = 24'b000000000000000111101010;
    16'b1111010010111101 : data_out = 24'b000000000000000111101010;
    16'b1111010010111110 : data_out = 24'b000000000000000111101011;
    16'b1111010010111111 : data_out = 24'b000000000000000111101011;
    16'b1111010011000000 : data_out = 24'b000000000000000111101011;
    16'b1111010011000001 : data_out = 24'b000000000000000111101100;
    16'b1111010011000010 : data_out = 24'b000000000000000111101100;
    16'b1111010011000011 : data_out = 24'b000000000000000111101101;
    16'b1111010011000100 : data_out = 24'b000000000000000111101101;
    16'b1111010011000101 : data_out = 24'b000000000000000111101110;
    16'b1111010011000110 : data_out = 24'b000000000000000111101110;
    16'b1111010011000111 : data_out = 24'b000000000000000111101111;
    16'b1111010011001000 : data_out = 24'b000000000000000111101111;
    16'b1111010011001001 : data_out = 24'b000000000000000111110000;
    16'b1111010011001010 : data_out = 24'b000000000000000111110000;
    16'b1111010011001011 : data_out = 24'b000000000000000111110001;
    16'b1111010011001100 : data_out = 24'b000000000000000111110001;
    16'b1111010011001101 : data_out = 24'b000000000000000111110010;
    16'b1111010011001110 : data_out = 24'b000000000000000111110010;
    16'b1111010011001111 : data_out = 24'b000000000000000111110011;
    16'b1111010011010000 : data_out = 24'b000000000000000111110011;
    16'b1111010011010001 : data_out = 24'b000000000000000111110100;
    16'b1111010011010010 : data_out = 24'b000000000000000111110100;
    16'b1111010011010011 : data_out = 24'b000000000000000111110101;
    16'b1111010011010100 : data_out = 24'b000000000000000111110101;
    16'b1111010011010101 : data_out = 24'b000000000000000111110110;
    16'b1111010011010110 : data_out = 24'b000000000000000111110110;
    16'b1111010011010111 : data_out = 24'b000000000000000111110111;
    16'b1111010011011000 : data_out = 24'b000000000000000111110111;
    16'b1111010011011001 : data_out = 24'b000000000000000111111000;
    16'b1111010011011010 : data_out = 24'b000000000000000111111000;
    16'b1111010011011011 : data_out = 24'b000000000000000111111001;
    16'b1111010011011100 : data_out = 24'b000000000000000111111001;
    16'b1111010011011101 : data_out = 24'b000000000000000111111010;
    16'b1111010011011110 : data_out = 24'b000000000000000111111010;
    16'b1111010011011111 : data_out = 24'b000000000000000111111011;
    16'b1111010011100000 : data_out = 24'b000000000000000111111011;
    16'b1111010011100001 : data_out = 24'b000000000000000111111100;
    16'b1111010011100010 : data_out = 24'b000000000000000111111100;
    16'b1111010011100011 : data_out = 24'b000000000000000111111101;
    16'b1111010011100100 : data_out = 24'b000000000000000111111101;
    16'b1111010011100101 : data_out = 24'b000000000000000111111110;
    16'b1111010011100110 : data_out = 24'b000000000000000111111110;
    16'b1111010011100111 : data_out = 24'b000000000000000111111111;
    16'b1111010011101000 : data_out = 24'b000000000000000111111111;
    16'b1111010011101001 : data_out = 24'b000000000000001000000000;
    16'b1111010011101010 : data_out = 24'b000000000000001000000000;
    16'b1111010011101011 : data_out = 24'b000000000000001000000001;
    16'b1111010011101100 : data_out = 24'b000000000000001000000001;
    16'b1111010011101101 : data_out = 24'b000000000000001000000010;
    16'b1111010011101110 : data_out = 24'b000000000000001000000010;
    16'b1111010011101111 : data_out = 24'b000000000000001000000011;
    16'b1111010011110000 : data_out = 24'b000000000000001000000011;
    16'b1111010011110001 : data_out = 24'b000000000000001000000100;
    16'b1111010011110010 : data_out = 24'b000000000000001000000100;
    16'b1111010011110011 : data_out = 24'b000000000000001000000101;
    16'b1111010011110100 : data_out = 24'b000000000000001000000101;
    16'b1111010011110101 : data_out = 24'b000000000000001000000110;
    16'b1111010011110110 : data_out = 24'b000000000000001000000110;
    16'b1111010011110111 : data_out = 24'b000000000000001000000111;
    16'b1111010011111000 : data_out = 24'b000000000000001000000111;
    16'b1111010011111001 : data_out = 24'b000000000000001000001000;
    16'b1111010011111010 : data_out = 24'b000000000000001000001000;
    16'b1111010011111011 : data_out = 24'b000000000000001000001001;
    16'b1111010011111100 : data_out = 24'b000000000000001000001001;
    16'b1111010011111101 : data_out = 24'b000000000000001000001010;
    16'b1111010011111110 : data_out = 24'b000000000000001000001010;
    16'b1111010011111111 : data_out = 24'b000000000000001000001011;
    16'b1111010100000000 : data_out = 24'b000000000000001000001011;
    16'b1111010100000001 : data_out = 24'b000000000000001000001100;
    16'b1111010100000010 : data_out = 24'b000000000000001000001100;
    16'b1111010100000011 : data_out = 24'b000000000000001000001101;
    16'b1111010100000100 : data_out = 24'b000000000000001000001101;
    16'b1111010100000101 : data_out = 24'b000000000000001000001110;
    16'b1111010100000110 : data_out = 24'b000000000000001000001110;
    16'b1111010100000111 : data_out = 24'b000000000000001000001111;
    16'b1111010100001000 : data_out = 24'b000000000000001000001111;
    16'b1111010100001001 : data_out = 24'b000000000000001000010000;
    16'b1111010100001010 : data_out = 24'b000000000000001000010000;
    16'b1111010100001011 : data_out = 24'b000000000000001000010001;
    16'b1111010100001100 : data_out = 24'b000000000000001000010001;
    16'b1111010100001101 : data_out = 24'b000000000000001000010010;
    16'b1111010100001110 : data_out = 24'b000000000000001000010010;
    16'b1111010100001111 : data_out = 24'b000000000000001000010011;
    16'b1111010100010000 : data_out = 24'b000000000000001000010011;
    16'b1111010100010001 : data_out = 24'b000000000000001000010100;
    16'b1111010100010010 : data_out = 24'b000000000000001000010100;
    16'b1111010100010011 : data_out = 24'b000000000000001000010101;
    16'b1111010100010100 : data_out = 24'b000000000000001000010110;
    16'b1111010100010101 : data_out = 24'b000000000000001000010110;
    16'b1111010100010110 : data_out = 24'b000000000000001000010111;
    16'b1111010100010111 : data_out = 24'b000000000000001000010111;
    16'b1111010100011000 : data_out = 24'b000000000000001000011000;
    16'b1111010100011001 : data_out = 24'b000000000000001000011000;
    16'b1111010100011010 : data_out = 24'b000000000000001000011001;
    16'b1111010100011011 : data_out = 24'b000000000000001000011001;
    16'b1111010100011100 : data_out = 24'b000000000000001000011010;
    16'b1111010100011101 : data_out = 24'b000000000000001000011010;
    16'b1111010100011110 : data_out = 24'b000000000000001000011011;
    16'b1111010100011111 : data_out = 24'b000000000000001000011011;
    16'b1111010100100000 : data_out = 24'b000000000000001000011100;
    16'b1111010100100001 : data_out = 24'b000000000000001000011100;
    16'b1111010100100010 : data_out = 24'b000000000000001000011101;
    16'b1111010100100011 : data_out = 24'b000000000000001000011101;
    16'b1111010100100100 : data_out = 24'b000000000000001000011110;
    16'b1111010100100101 : data_out = 24'b000000000000001000011110;
    16'b1111010100100110 : data_out = 24'b000000000000001000011111;
    16'b1111010100100111 : data_out = 24'b000000000000001000100000;
    16'b1111010100101000 : data_out = 24'b000000000000001000100000;
    16'b1111010100101001 : data_out = 24'b000000000000001000100001;
    16'b1111010100101010 : data_out = 24'b000000000000001000100001;
    16'b1111010100101011 : data_out = 24'b000000000000001000100010;
    16'b1111010100101100 : data_out = 24'b000000000000001000100010;
    16'b1111010100101101 : data_out = 24'b000000000000001000100011;
    16'b1111010100101110 : data_out = 24'b000000000000001000100011;
    16'b1111010100101111 : data_out = 24'b000000000000001000100100;
    16'b1111010100110000 : data_out = 24'b000000000000001000100100;
    16'b1111010100110001 : data_out = 24'b000000000000001000100101;
    16'b1111010100110010 : data_out = 24'b000000000000001000100101;
    16'b1111010100110011 : data_out = 24'b000000000000001000100110;
    16'b1111010100110100 : data_out = 24'b000000000000001000100110;
    16'b1111010100110101 : data_out = 24'b000000000000001000100111;
    16'b1111010100110110 : data_out = 24'b000000000000001000101000;
    16'b1111010100110111 : data_out = 24'b000000000000001000101000;
    16'b1111010100111000 : data_out = 24'b000000000000001000101001;
    16'b1111010100111001 : data_out = 24'b000000000000001000101001;
    16'b1111010100111010 : data_out = 24'b000000000000001000101010;
    16'b1111010100111011 : data_out = 24'b000000000000001000101010;
    16'b1111010100111100 : data_out = 24'b000000000000001000101011;
    16'b1111010100111101 : data_out = 24'b000000000000001000101011;
    16'b1111010100111110 : data_out = 24'b000000000000001000101100;
    16'b1111010100111111 : data_out = 24'b000000000000001000101100;
    16'b1111010101000000 : data_out = 24'b000000000000001000101101;
    16'b1111010101000001 : data_out = 24'b000000000000001000101110;
    16'b1111010101000010 : data_out = 24'b000000000000001000101110;
    16'b1111010101000011 : data_out = 24'b000000000000001000101111;
    16'b1111010101000100 : data_out = 24'b000000000000001000101111;
    16'b1111010101000101 : data_out = 24'b000000000000001000110000;
    16'b1111010101000110 : data_out = 24'b000000000000001000110000;
    16'b1111010101000111 : data_out = 24'b000000000000001000110001;
    16'b1111010101001000 : data_out = 24'b000000000000001000110001;
    16'b1111010101001001 : data_out = 24'b000000000000001000110010;
    16'b1111010101001010 : data_out = 24'b000000000000001000110010;
    16'b1111010101001011 : data_out = 24'b000000000000001000110011;
    16'b1111010101001100 : data_out = 24'b000000000000001000110100;
    16'b1111010101001101 : data_out = 24'b000000000000001000110100;
    16'b1111010101001110 : data_out = 24'b000000000000001000110101;
    16'b1111010101001111 : data_out = 24'b000000000000001000110101;
    16'b1111010101010000 : data_out = 24'b000000000000001000110110;
    16'b1111010101010001 : data_out = 24'b000000000000001000110110;
    16'b1111010101010010 : data_out = 24'b000000000000001000110111;
    16'b1111010101010011 : data_out = 24'b000000000000001000110111;
    16'b1111010101010100 : data_out = 24'b000000000000001000111000;
    16'b1111010101010101 : data_out = 24'b000000000000001000111001;
    16'b1111010101010110 : data_out = 24'b000000000000001000111001;
    16'b1111010101010111 : data_out = 24'b000000000000001000111010;
    16'b1111010101011000 : data_out = 24'b000000000000001000111010;
    16'b1111010101011001 : data_out = 24'b000000000000001000111011;
    16'b1111010101011010 : data_out = 24'b000000000000001000111011;
    16'b1111010101011011 : data_out = 24'b000000000000001000111100;
    16'b1111010101011100 : data_out = 24'b000000000000001000111100;
    16'b1111010101011101 : data_out = 24'b000000000000001000111101;
    16'b1111010101011110 : data_out = 24'b000000000000001000111110;
    16'b1111010101011111 : data_out = 24'b000000000000001000111110;
    16'b1111010101100000 : data_out = 24'b000000000000001000111111;
    16'b1111010101100001 : data_out = 24'b000000000000001000111111;
    16'b1111010101100010 : data_out = 24'b000000000000001001000000;
    16'b1111010101100011 : data_out = 24'b000000000000001001000000;
    16'b1111010101100100 : data_out = 24'b000000000000001001000001;
    16'b1111010101100101 : data_out = 24'b000000000000001001000001;
    16'b1111010101100110 : data_out = 24'b000000000000001001000010;
    16'b1111010101100111 : data_out = 24'b000000000000001001000011;
    16'b1111010101101000 : data_out = 24'b000000000000001001000011;
    16'b1111010101101001 : data_out = 24'b000000000000001001000100;
    16'b1111010101101010 : data_out = 24'b000000000000001001000100;
    16'b1111010101101011 : data_out = 24'b000000000000001001000101;
    16'b1111010101101100 : data_out = 24'b000000000000001001000101;
    16'b1111010101101101 : data_out = 24'b000000000000001001000110;
    16'b1111010101101110 : data_out = 24'b000000000000001001000111;
    16'b1111010101101111 : data_out = 24'b000000000000001001000111;
    16'b1111010101110000 : data_out = 24'b000000000000001001001000;
    16'b1111010101110001 : data_out = 24'b000000000000001001001000;
    16'b1111010101110010 : data_out = 24'b000000000000001001001001;
    16'b1111010101110011 : data_out = 24'b000000000000001001001001;
    16'b1111010101110100 : data_out = 24'b000000000000001001001010;
    16'b1111010101110101 : data_out = 24'b000000000000001001001011;
    16'b1111010101110110 : data_out = 24'b000000000000001001001011;
    16'b1111010101110111 : data_out = 24'b000000000000001001001100;
    16'b1111010101111000 : data_out = 24'b000000000000001001001100;
    16'b1111010101111001 : data_out = 24'b000000000000001001001101;
    16'b1111010101111010 : data_out = 24'b000000000000001001001101;
    16'b1111010101111011 : data_out = 24'b000000000000001001001110;
    16'b1111010101111100 : data_out = 24'b000000000000001001001111;
    16'b1111010101111101 : data_out = 24'b000000000000001001001111;
    16'b1111010101111110 : data_out = 24'b000000000000001001010000;
    16'b1111010101111111 : data_out = 24'b000000000000001001010000;
    16'b1111010110000000 : data_out = 24'b000000000000001001010001;
    16'b1111010110000001 : data_out = 24'b000000000000001001010010;
    16'b1111010110000010 : data_out = 24'b000000000000001001010010;
    16'b1111010110000011 : data_out = 24'b000000000000001001010011;
    16'b1111010110000100 : data_out = 24'b000000000000001001010011;
    16'b1111010110000101 : data_out = 24'b000000000000001001010100;
    16'b1111010110000110 : data_out = 24'b000000000000001001010100;
    16'b1111010110000111 : data_out = 24'b000000000000001001010101;
    16'b1111010110001000 : data_out = 24'b000000000000001001010110;
    16'b1111010110001001 : data_out = 24'b000000000000001001010110;
    16'b1111010110001010 : data_out = 24'b000000000000001001010111;
    16'b1111010110001011 : data_out = 24'b000000000000001001010111;
    16'b1111010110001100 : data_out = 24'b000000000000001001011000;
    16'b1111010110001101 : data_out = 24'b000000000000001001011001;
    16'b1111010110001110 : data_out = 24'b000000000000001001011001;
    16'b1111010110001111 : data_out = 24'b000000000000001001011010;
    16'b1111010110010000 : data_out = 24'b000000000000001001011010;
    16'b1111010110010001 : data_out = 24'b000000000000001001011011;
    16'b1111010110010010 : data_out = 24'b000000000000001001011011;
    16'b1111010110010011 : data_out = 24'b000000000000001001011100;
    16'b1111010110010100 : data_out = 24'b000000000000001001011101;
    16'b1111010110010101 : data_out = 24'b000000000000001001011101;
    16'b1111010110010110 : data_out = 24'b000000000000001001011110;
    16'b1111010110010111 : data_out = 24'b000000000000001001011110;
    16'b1111010110011000 : data_out = 24'b000000000000001001011111;
    16'b1111010110011001 : data_out = 24'b000000000000001001100000;
    16'b1111010110011010 : data_out = 24'b000000000000001001100000;
    16'b1111010110011011 : data_out = 24'b000000000000001001100001;
    16'b1111010110011100 : data_out = 24'b000000000000001001100001;
    16'b1111010110011101 : data_out = 24'b000000000000001001100010;
    16'b1111010110011110 : data_out = 24'b000000000000001001100011;
    16'b1111010110011111 : data_out = 24'b000000000000001001100011;
    16'b1111010110100000 : data_out = 24'b000000000000001001100100;
    16'b1111010110100001 : data_out = 24'b000000000000001001100100;
    16'b1111010110100010 : data_out = 24'b000000000000001001100101;
    16'b1111010110100011 : data_out = 24'b000000000000001001100110;
    16'b1111010110100100 : data_out = 24'b000000000000001001100110;
    16'b1111010110100101 : data_out = 24'b000000000000001001100111;
    16'b1111010110100110 : data_out = 24'b000000000000001001100111;
    16'b1111010110100111 : data_out = 24'b000000000000001001101000;
    16'b1111010110101000 : data_out = 24'b000000000000001001101001;
    16'b1111010110101001 : data_out = 24'b000000000000001001101001;
    16'b1111010110101010 : data_out = 24'b000000000000001001101010;
    16'b1111010110101011 : data_out = 24'b000000000000001001101010;
    16'b1111010110101100 : data_out = 24'b000000000000001001101011;
    16'b1111010110101101 : data_out = 24'b000000000000001001101100;
    16'b1111010110101110 : data_out = 24'b000000000000001001101100;
    16'b1111010110101111 : data_out = 24'b000000000000001001101101;
    16'b1111010110110000 : data_out = 24'b000000000000001001101101;
    16'b1111010110110001 : data_out = 24'b000000000000001001101110;
    16'b1111010110110010 : data_out = 24'b000000000000001001101111;
    16'b1111010110110011 : data_out = 24'b000000000000001001101111;
    16'b1111010110110100 : data_out = 24'b000000000000001001110000;
    16'b1111010110110101 : data_out = 24'b000000000000001001110000;
    16'b1111010110110110 : data_out = 24'b000000000000001001110001;
    16'b1111010110110111 : data_out = 24'b000000000000001001110010;
    16'b1111010110111000 : data_out = 24'b000000000000001001110010;
    16'b1111010110111001 : data_out = 24'b000000000000001001110011;
    16'b1111010110111010 : data_out = 24'b000000000000001001110100;
    16'b1111010110111011 : data_out = 24'b000000000000001001110100;
    16'b1111010110111100 : data_out = 24'b000000000000001001110101;
    16'b1111010110111101 : data_out = 24'b000000000000001001110101;
    16'b1111010110111110 : data_out = 24'b000000000000001001110110;
    16'b1111010110111111 : data_out = 24'b000000000000001001110111;
    16'b1111010111000000 : data_out = 24'b000000000000001001110111;
    16'b1111010111000001 : data_out = 24'b000000000000001001111000;
    16'b1111010111000010 : data_out = 24'b000000000000001001111000;
    16'b1111010111000011 : data_out = 24'b000000000000001001111001;
    16'b1111010111000100 : data_out = 24'b000000000000001001111010;
    16'b1111010111000101 : data_out = 24'b000000000000001001111010;
    16'b1111010111000110 : data_out = 24'b000000000000001001111011;
    16'b1111010111000111 : data_out = 24'b000000000000001001111100;
    16'b1111010111001000 : data_out = 24'b000000000000001001111100;
    16'b1111010111001001 : data_out = 24'b000000000000001001111101;
    16'b1111010111001010 : data_out = 24'b000000000000001001111101;
    16'b1111010111001011 : data_out = 24'b000000000000001001111110;
    16'b1111010111001100 : data_out = 24'b000000000000001001111111;
    16'b1111010111001101 : data_out = 24'b000000000000001001111111;
    16'b1111010111001110 : data_out = 24'b000000000000001010000000;
    16'b1111010111001111 : data_out = 24'b000000000000001010000001;
    16'b1111010111010000 : data_out = 24'b000000000000001010000001;
    16'b1111010111010001 : data_out = 24'b000000000000001010000010;
    16'b1111010111010010 : data_out = 24'b000000000000001010000010;
    16'b1111010111010011 : data_out = 24'b000000000000001010000011;
    16'b1111010111010100 : data_out = 24'b000000000000001010000100;
    16'b1111010111010101 : data_out = 24'b000000000000001010000100;
    16'b1111010111010110 : data_out = 24'b000000000000001010000101;
    16'b1111010111010111 : data_out = 24'b000000000000001010000110;
    16'b1111010111011000 : data_out = 24'b000000000000001010000110;
    16'b1111010111011001 : data_out = 24'b000000000000001010000111;
    16'b1111010111011010 : data_out = 24'b000000000000001010000111;
    16'b1111010111011011 : data_out = 24'b000000000000001010001000;
    16'b1111010111011100 : data_out = 24'b000000000000001010001001;
    16'b1111010111011101 : data_out = 24'b000000000000001010001001;
    16'b1111010111011110 : data_out = 24'b000000000000001010001010;
    16'b1111010111011111 : data_out = 24'b000000000000001010001011;
    16'b1111010111100000 : data_out = 24'b000000000000001010001011;
    16'b1111010111100001 : data_out = 24'b000000000000001010001100;
    16'b1111010111100010 : data_out = 24'b000000000000001010001101;
    16'b1111010111100011 : data_out = 24'b000000000000001010001101;
    16'b1111010111100100 : data_out = 24'b000000000000001010001110;
    16'b1111010111100101 : data_out = 24'b000000000000001010001110;
    16'b1111010111100110 : data_out = 24'b000000000000001010001111;
    16'b1111010111100111 : data_out = 24'b000000000000001010010000;
    16'b1111010111101000 : data_out = 24'b000000000000001010010000;
    16'b1111010111101001 : data_out = 24'b000000000000001010010001;
    16'b1111010111101010 : data_out = 24'b000000000000001010010010;
    16'b1111010111101011 : data_out = 24'b000000000000001010010010;
    16'b1111010111101100 : data_out = 24'b000000000000001010010011;
    16'b1111010111101101 : data_out = 24'b000000000000001010010100;
    16'b1111010111101110 : data_out = 24'b000000000000001010010100;
    16'b1111010111101111 : data_out = 24'b000000000000001010010101;
    16'b1111010111110000 : data_out = 24'b000000000000001010010110;
    16'b1111010111110001 : data_out = 24'b000000000000001010010110;
    16'b1111010111110010 : data_out = 24'b000000000000001010010111;
    16'b1111010111110011 : data_out = 24'b000000000000001010010111;
    16'b1111010111110100 : data_out = 24'b000000000000001010011000;
    16'b1111010111110101 : data_out = 24'b000000000000001010011001;
    16'b1111010111110110 : data_out = 24'b000000000000001010011001;
    16'b1111010111110111 : data_out = 24'b000000000000001010011010;
    16'b1111010111111000 : data_out = 24'b000000000000001010011011;
    16'b1111010111111001 : data_out = 24'b000000000000001010011011;
    16'b1111010111111010 : data_out = 24'b000000000000001010011100;
    16'b1111010111111011 : data_out = 24'b000000000000001010011101;
    16'b1111010111111100 : data_out = 24'b000000000000001010011101;
    16'b1111010111111101 : data_out = 24'b000000000000001010011110;
    16'b1111010111111110 : data_out = 24'b000000000000001010011111;
    16'b1111010111111111 : data_out = 24'b000000000000001010011111;
    16'b1111011000000000 : data_out = 24'b000000000000001010100000;
    16'b1111011000000001 : data_out = 24'b000000000000001010100001;
    16'b1111011000000010 : data_out = 24'b000000000000001010100001;
    16'b1111011000000011 : data_out = 24'b000000000000001010100010;
    16'b1111011000000100 : data_out = 24'b000000000000001010100011;
    16'b1111011000000101 : data_out = 24'b000000000000001010100011;
    16'b1111011000000110 : data_out = 24'b000000000000001010100100;
    16'b1111011000000111 : data_out = 24'b000000000000001010100101;
    16'b1111011000001000 : data_out = 24'b000000000000001010100101;
    16'b1111011000001001 : data_out = 24'b000000000000001010100110;
    16'b1111011000001010 : data_out = 24'b000000000000001010100111;
    16'b1111011000001011 : data_out = 24'b000000000000001010100111;
    16'b1111011000001100 : data_out = 24'b000000000000001010101000;
    16'b1111011000001101 : data_out = 24'b000000000000001010101001;
    16'b1111011000001110 : data_out = 24'b000000000000001010101001;
    16'b1111011000001111 : data_out = 24'b000000000000001010101010;
    16'b1111011000010000 : data_out = 24'b000000000000001010101011;
    16'b1111011000010001 : data_out = 24'b000000000000001010101011;
    16'b1111011000010010 : data_out = 24'b000000000000001010101100;
    16'b1111011000010011 : data_out = 24'b000000000000001010101101;
    16'b1111011000010100 : data_out = 24'b000000000000001010101101;
    16'b1111011000010101 : data_out = 24'b000000000000001010101110;
    16'b1111011000010110 : data_out = 24'b000000000000001010101111;
    16'b1111011000010111 : data_out = 24'b000000000000001010101111;
    16'b1111011000011000 : data_out = 24'b000000000000001010110000;
    16'b1111011000011001 : data_out = 24'b000000000000001010110001;
    16'b1111011000011010 : data_out = 24'b000000000000001010110001;
    16'b1111011000011011 : data_out = 24'b000000000000001010110010;
    16'b1111011000011100 : data_out = 24'b000000000000001010110011;
    16'b1111011000011101 : data_out = 24'b000000000000001010110011;
    16'b1111011000011110 : data_out = 24'b000000000000001010110100;
    16'b1111011000011111 : data_out = 24'b000000000000001010110101;
    16'b1111011000100000 : data_out = 24'b000000000000001010110101;
    16'b1111011000100001 : data_out = 24'b000000000000001010110110;
    16'b1111011000100010 : data_out = 24'b000000000000001010110111;
    16'b1111011000100011 : data_out = 24'b000000000000001010110111;
    16'b1111011000100100 : data_out = 24'b000000000000001010111000;
    16'b1111011000100101 : data_out = 24'b000000000000001010111001;
    16'b1111011000100110 : data_out = 24'b000000000000001010111001;
    16'b1111011000100111 : data_out = 24'b000000000000001010111010;
    16'b1111011000101000 : data_out = 24'b000000000000001010111011;
    16'b1111011000101001 : data_out = 24'b000000000000001010111011;
    16'b1111011000101010 : data_out = 24'b000000000000001010111100;
    16'b1111011000101011 : data_out = 24'b000000000000001010111101;
    16'b1111011000101100 : data_out = 24'b000000000000001010111101;
    16'b1111011000101101 : data_out = 24'b000000000000001010111110;
    16'b1111011000101110 : data_out = 24'b000000000000001010111111;
    16'b1111011000101111 : data_out = 24'b000000000000001011000000;
    16'b1111011000110000 : data_out = 24'b000000000000001011000000;
    16'b1111011000110001 : data_out = 24'b000000000000001011000001;
    16'b1111011000110010 : data_out = 24'b000000000000001011000010;
    16'b1111011000110011 : data_out = 24'b000000000000001011000010;
    16'b1111011000110100 : data_out = 24'b000000000000001011000011;
    16'b1111011000110101 : data_out = 24'b000000000000001011000100;
    16'b1111011000110110 : data_out = 24'b000000000000001011000100;
    16'b1111011000110111 : data_out = 24'b000000000000001011000101;
    16'b1111011000111000 : data_out = 24'b000000000000001011000110;
    16'b1111011000111001 : data_out = 24'b000000000000001011000110;
    16'b1111011000111010 : data_out = 24'b000000000000001011000111;
    16'b1111011000111011 : data_out = 24'b000000000000001011001000;
    16'b1111011000111100 : data_out = 24'b000000000000001011001001;
    16'b1111011000111101 : data_out = 24'b000000000000001011001001;
    16'b1111011000111110 : data_out = 24'b000000000000001011001010;
    16'b1111011000111111 : data_out = 24'b000000000000001011001011;
    16'b1111011001000000 : data_out = 24'b000000000000001011001011;
    16'b1111011001000001 : data_out = 24'b000000000000001011001100;
    16'b1111011001000010 : data_out = 24'b000000000000001011001101;
    16'b1111011001000011 : data_out = 24'b000000000000001011001101;
    16'b1111011001000100 : data_out = 24'b000000000000001011001110;
    16'b1111011001000101 : data_out = 24'b000000000000001011001111;
    16'b1111011001000110 : data_out = 24'b000000000000001011010000;
    16'b1111011001000111 : data_out = 24'b000000000000001011010000;
    16'b1111011001001000 : data_out = 24'b000000000000001011010001;
    16'b1111011001001001 : data_out = 24'b000000000000001011010010;
    16'b1111011001001010 : data_out = 24'b000000000000001011010010;
    16'b1111011001001011 : data_out = 24'b000000000000001011010011;
    16'b1111011001001100 : data_out = 24'b000000000000001011010100;
    16'b1111011001001101 : data_out = 24'b000000000000001011010100;
    16'b1111011001001110 : data_out = 24'b000000000000001011010101;
    16'b1111011001001111 : data_out = 24'b000000000000001011010110;
    16'b1111011001010000 : data_out = 24'b000000000000001011010111;
    16'b1111011001010001 : data_out = 24'b000000000000001011010111;
    16'b1111011001010010 : data_out = 24'b000000000000001011011000;
    16'b1111011001010011 : data_out = 24'b000000000000001011011001;
    16'b1111011001010100 : data_out = 24'b000000000000001011011001;
    16'b1111011001010101 : data_out = 24'b000000000000001011011010;
    16'b1111011001010110 : data_out = 24'b000000000000001011011011;
    16'b1111011001010111 : data_out = 24'b000000000000001011011100;
    16'b1111011001011000 : data_out = 24'b000000000000001011011100;
    16'b1111011001011001 : data_out = 24'b000000000000001011011101;
    16'b1111011001011010 : data_out = 24'b000000000000001011011110;
    16'b1111011001011011 : data_out = 24'b000000000000001011011110;
    16'b1111011001011100 : data_out = 24'b000000000000001011011111;
    16'b1111011001011101 : data_out = 24'b000000000000001011100000;
    16'b1111011001011110 : data_out = 24'b000000000000001011100001;
    16'b1111011001011111 : data_out = 24'b000000000000001011100001;
    16'b1111011001100000 : data_out = 24'b000000000000001011100010;
    16'b1111011001100001 : data_out = 24'b000000000000001011100011;
    16'b1111011001100010 : data_out = 24'b000000000000001011100011;
    16'b1111011001100011 : data_out = 24'b000000000000001011100100;
    16'b1111011001100100 : data_out = 24'b000000000000001011100101;
    16'b1111011001100101 : data_out = 24'b000000000000001011100110;
    16'b1111011001100110 : data_out = 24'b000000000000001011100110;
    16'b1111011001100111 : data_out = 24'b000000000000001011100111;
    16'b1111011001101000 : data_out = 24'b000000000000001011101000;
    16'b1111011001101001 : data_out = 24'b000000000000001011101001;
    16'b1111011001101010 : data_out = 24'b000000000000001011101001;
    16'b1111011001101011 : data_out = 24'b000000000000001011101010;
    16'b1111011001101100 : data_out = 24'b000000000000001011101011;
    16'b1111011001101101 : data_out = 24'b000000000000001011101011;
    16'b1111011001101110 : data_out = 24'b000000000000001011101100;
    16'b1111011001101111 : data_out = 24'b000000000000001011101101;
    16'b1111011001110000 : data_out = 24'b000000000000001011101110;
    16'b1111011001110001 : data_out = 24'b000000000000001011101110;
    16'b1111011001110010 : data_out = 24'b000000000000001011101111;
    16'b1111011001110011 : data_out = 24'b000000000000001011110000;
    16'b1111011001110100 : data_out = 24'b000000000000001011110001;
    16'b1111011001110101 : data_out = 24'b000000000000001011110001;
    16'b1111011001110110 : data_out = 24'b000000000000001011110010;
    16'b1111011001110111 : data_out = 24'b000000000000001011110011;
    16'b1111011001111000 : data_out = 24'b000000000000001011110100;
    16'b1111011001111001 : data_out = 24'b000000000000001011110100;
    16'b1111011001111010 : data_out = 24'b000000000000001011110101;
    16'b1111011001111011 : data_out = 24'b000000000000001011110110;
    16'b1111011001111100 : data_out = 24'b000000000000001011110111;
    16'b1111011001111101 : data_out = 24'b000000000000001011110111;
    16'b1111011001111110 : data_out = 24'b000000000000001011111000;
    16'b1111011001111111 : data_out = 24'b000000000000001011111001;
    16'b1111011010000000 : data_out = 24'b000000000000001011111001;
    16'b1111011010000001 : data_out = 24'b000000000000001011111010;
    16'b1111011010000010 : data_out = 24'b000000000000001011111011;
    16'b1111011010000011 : data_out = 24'b000000000000001011111100;
    16'b1111011010000100 : data_out = 24'b000000000000001011111100;
    16'b1111011010000101 : data_out = 24'b000000000000001011111101;
    16'b1111011010000110 : data_out = 24'b000000000000001011111110;
    16'b1111011010000111 : data_out = 24'b000000000000001011111111;
    16'b1111011010001000 : data_out = 24'b000000000000001011111111;
    16'b1111011010001001 : data_out = 24'b000000000000001100000000;
    16'b1111011010001010 : data_out = 24'b000000000000001100000001;
    16'b1111011010001011 : data_out = 24'b000000000000001100000010;
    16'b1111011010001100 : data_out = 24'b000000000000001100000010;
    16'b1111011010001101 : data_out = 24'b000000000000001100000011;
    16'b1111011010001110 : data_out = 24'b000000000000001100000100;
    16'b1111011010001111 : data_out = 24'b000000000000001100000101;
    16'b1111011010010000 : data_out = 24'b000000000000001100000101;
    16'b1111011010010001 : data_out = 24'b000000000000001100000110;
    16'b1111011010010010 : data_out = 24'b000000000000001100000111;
    16'b1111011010010011 : data_out = 24'b000000000000001100001000;
    16'b1111011010010100 : data_out = 24'b000000000000001100001001;
    16'b1111011010010101 : data_out = 24'b000000000000001100001001;
    16'b1111011010010110 : data_out = 24'b000000000000001100001010;
    16'b1111011010010111 : data_out = 24'b000000000000001100001011;
    16'b1111011010011000 : data_out = 24'b000000000000001100001100;
    16'b1111011010011001 : data_out = 24'b000000000000001100001100;
    16'b1111011010011010 : data_out = 24'b000000000000001100001101;
    16'b1111011010011011 : data_out = 24'b000000000000001100001110;
    16'b1111011010011100 : data_out = 24'b000000000000001100001111;
    16'b1111011010011101 : data_out = 24'b000000000000001100001111;
    16'b1111011010011110 : data_out = 24'b000000000000001100010000;
    16'b1111011010011111 : data_out = 24'b000000000000001100010001;
    16'b1111011010100000 : data_out = 24'b000000000000001100010010;
    16'b1111011010100001 : data_out = 24'b000000000000001100010010;
    16'b1111011010100010 : data_out = 24'b000000000000001100010011;
    16'b1111011010100011 : data_out = 24'b000000000000001100010100;
    16'b1111011010100100 : data_out = 24'b000000000000001100010101;
    16'b1111011010100101 : data_out = 24'b000000000000001100010110;
    16'b1111011010100110 : data_out = 24'b000000000000001100010110;
    16'b1111011010100111 : data_out = 24'b000000000000001100010111;
    16'b1111011010101000 : data_out = 24'b000000000000001100011000;
    16'b1111011010101001 : data_out = 24'b000000000000001100011001;
    16'b1111011010101010 : data_out = 24'b000000000000001100011001;
    16'b1111011010101011 : data_out = 24'b000000000000001100011010;
    16'b1111011010101100 : data_out = 24'b000000000000001100011011;
    16'b1111011010101101 : data_out = 24'b000000000000001100011100;
    16'b1111011010101110 : data_out = 24'b000000000000001100011100;
    16'b1111011010101111 : data_out = 24'b000000000000001100011101;
    16'b1111011010110000 : data_out = 24'b000000000000001100011110;
    16'b1111011010110001 : data_out = 24'b000000000000001100011111;
    16'b1111011010110010 : data_out = 24'b000000000000001100100000;
    16'b1111011010110011 : data_out = 24'b000000000000001100100000;
    16'b1111011010110100 : data_out = 24'b000000000000001100100001;
    16'b1111011010110101 : data_out = 24'b000000000000001100100010;
    16'b1111011010110110 : data_out = 24'b000000000000001100100011;
    16'b1111011010110111 : data_out = 24'b000000000000001100100100;
    16'b1111011010111000 : data_out = 24'b000000000000001100100100;
    16'b1111011010111001 : data_out = 24'b000000000000001100100101;
    16'b1111011010111010 : data_out = 24'b000000000000001100100110;
    16'b1111011010111011 : data_out = 24'b000000000000001100100111;
    16'b1111011010111100 : data_out = 24'b000000000000001100100111;
    16'b1111011010111101 : data_out = 24'b000000000000001100101000;
    16'b1111011010111110 : data_out = 24'b000000000000001100101001;
    16'b1111011010111111 : data_out = 24'b000000000000001100101010;
    16'b1111011011000000 : data_out = 24'b000000000000001100101011;
    16'b1111011011000001 : data_out = 24'b000000000000001100101011;
    16'b1111011011000010 : data_out = 24'b000000000000001100101100;
    16'b1111011011000011 : data_out = 24'b000000000000001100101101;
    16'b1111011011000100 : data_out = 24'b000000000000001100101110;
    16'b1111011011000101 : data_out = 24'b000000000000001100101111;
    16'b1111011011000110 : data_out = 24'b000000000000001100101111;
    16'b1111011011000111 : data_out = 24'b000000000000001100110000;
    16'b1111011011001000 : data_out = 24'b000000000000001100110001;
    16'b1111011011001001 : data_out = 24'b000000000000001100110010;
    16'b1111011011001010 : data_out = 24'b000000000000001100110011;
    16'b1111011011001011 : data_out = 24'b000000000000001100110011;
    16'b1111011011001100 : data_out = 24'b000000000000001100110100;
    16'b1111011011001101 : data_out = 24'b000000000000001100110101;
    16'b1111011011001110 : data_out = 24'b000000000000001100110110;
    16'b1111011011001111 : data_out = 24'b000000000000001100110111;
    16'b1111011011010000 : data_out = 24'b000000000000001100110111;
    16'b1111011011010001 : data_out = 24'b000000000000001100111000;
    16'b1111011011010010 : data_out = 24'b000000000000001100111001;
    16'b1111011011010011 : data_out = 24'b000000000000001100111010;
    16'b1111011011010100 : data_out = 24'b000000000000001100111011;
    16'b1111011011010101 : data_out = 24'b000000000000001100111011;
    16'b1111011011010110 : data_out = 24'b000000000000001100111100;
    16'b1111011011010111 : data_out = 24'b000000000000001100111101;
    16'b1111011011011000 : data_out = 24'b000000000000001100111110;
    16'b1111011011011001 : data_out = 24'b000000000000001100111111;
    16'b1111011011011010 : data_out = 24'b000000000000001100111111;
    16'b1111011011011011 : data_out = 24'b000000000000001101000000;
    16'b1111011011011100 : data_out = 24'b000000000000001101000001;
    16'b1111011011011101 : data_out = 24'b000000000000001101000010;
    16'b1111011011011110 : data_out = 24'b000000000000001101000011;
    16'b1111011011011111 : data_out = 24'b000000000000001101000100;
    16'b1111011011100000 : data_out = 24'b000000000000001101000100;
    16'b1111011011100001 : data_out = 24'b000000000000001101000101;
    16'b1111011011100010 : data_out = 24'b000000000000001101000110;
    16'b1111011011100011 : data_out = 24'b000000000000001101000111;
    16'b1111011011100100 : data_out = 24'b000000000000001101001000;
    16'b1111011011100101 : data_out = 24'b000000000000001101001000;
    16'b1111011011100110 : data_out = 24'b000000000000001101001001;
    16'b1111011011100111 : data_out = 24'b000000000000001101001010;
    16'b1111011011101000 : data_out = 24'b000000000000001101001011;
    16'b1111011011101001 : data_out = 24'b000000000000001101001100;
    16'b1111011011101010 : data_out = 24'b000000000000001101001101;
    16'b1111011011101011 : data_out = 24'b000000000000001101001101;
    16'b1111011011101100 : data_out = 24'b000000000000001101001110;
    16'b1111011011101101 : data_out = 24'b000000000000001101001111;
    16'b1111011011101110 : data_out = 24'b000000000000001101010000;
    16'b1111011011101111 : data_out = 24'b000000000000001101010001;
    16'b1111011011110000 : data_out = 24'b000000000000001101010010;
    16'b1111011011110001 : data_out = 24'b000000000000001101010010;
    16'b1111011011110010 : data_out = 24'b000000000000001101010011;
    16'b1111011011110011 : data_out = 24'b000000000000001101010100;
    16'b1111011011110100 : data_out = 24'b000000000000001101010101;
    16'b1111011011110101 : data_out = 24'b000000000000001101010110;
    16'b1111011011110110 : data_out = 24'b000000000000001101010111;
    16'b1111011011110111 : data_out = 24'b000000000000001101010111;
    16'b1111011011111000 : data_out = 24'b000000000000001101011000;
    16'b1111011011111001 : data_out = 24'b000000000000001101011001;
    16'b1111011011111010 : data_out = 24'b000000000000001101011010;
    16'b1111011011111011 : data_out = 24'b000000000000001101011011;
    16'b1111011011111100 : data_out = 24'b000000000000001101011100;
    16'b1111011011111101 : data_out = 24'b000000000000001101011100;
    16'b1111011011111110 : data_out = 24'b000000000000001101011101;
    16'b1111011011111111 : data_out = 24'b000000000000001101011110;
    16'b1111011100000000 : data_out = 24'b000000000000001101011111;
    16'b1111011100000001 : data_out = 24'b000000000000001101100000;
    16'b1111011100000010 : data_out = 24'b000000000000001101100001;
    16'b1111011100000011 : data_out = 24'b000000000000001101100001;
    16'b1111011100000100 : data_out = 24'b000000000000001101100010;
    16'b1111011100000101 : data_out = 24'b000000000000001101100011;
    16'b1111011100000110 : data_out = 24'b000000000000001101100100;
    16'b1111011100000111 : data_out = 24'b000000000000001101100101;
    16'b1111011100001000 : data_out = 24'b000000000000001101100110;
    16'b1111011100001001 : data_out = 24'b000000000000001101100111;
    16'b1111011100001010 : data_out = 24'b000000000000001101100111;
    16'b1111011100001011 : data_out = 24'b000000000000001101101000;
    16'b1111011100001100 : data_out = 24'b000000000000001101101001;
    16'b1111011100001101 : data_out = 24'b000000000000001101101010;
    16'b1111011100001110 : data_out = 24'b000000000000001101101011;
    16'b1111011100001111 : data_out = 24'b000000000000001101101100;
    16'b1111011100010000 : data_out = 24'b000000000000001101101101;
    16'b1111011100010001 : data_out = 24'b000000000000001101101101;
    16'b1111011100010010 : data_out = 24'b000000000000001101101110;
    16'b1111011100010011 : data_out = 24'b000000000000001101101111;
    16'b1111011100010100 : data_out = 24'b000000000000001101110000;
    16'b1111011100010101 : data_out = 24'b000000000000001101110001;
    16'b1111011100010110 : data_out = 24'b000000000000001101110010;
    16'b1111011100010111 : data_out = 24'b000000000000001101110011;
    16'b1111011100011000 : data_out = 24'b000000000000001101110011;
    16'b1111011100011001 : data_out = 24'b000000000000001101110100;
    16'b1111011100011010 : data_out = 24'b000000000000001101110101;
    16'b1111011100011011 : data_out = 24'b000000000000001101110110;
    16'b1111011100011100 : data_out = 24'b000000000000001101110111;
    16'b1111011100011101 : data_out = 24'b000000000000001101111000;
    16'b1111011100011110 : data_out = 24'b000000000000001101111001;
    16'b1111011100011111 : data_out = 24'b000000000000001101111001;
    16'b1111011100100000 : data_out = 24'b000000000000001101111010;
    16'b1111011100100001 : data_out = 24'b000000000000001101111011;
    16'b1111011100100010 : data_out = 24'b000000000000001101111100;
    16'b1111011100100011 : data_out = 24'b000000000000001101111101;
    16'b1111011100100100 : data_out = 24'b000000000000001101111110;
    16'b1111011100100101 : data_out = 24'b000000000000001101111111;
    16'b1111011100100110 : data_out = 24'b000000000000001110000000;
    16'b1111011100100111 : data_out = 24'b000000000000001110000000;
    16'b1111011100101000 : data_out = 24'b000000000000001110000001;
    16'b1111011100101001 : data_out = 24'b000000000000001110000010;
    16'b1111011100101010 : data_out = 24'b000000000000001110000011;
    16'b1111011100101011 : data_out = 24'b000000000000001110000100;
    16'b1111011100101100 : data_out = 24'b000000000000001110000101;
    16'b1111011100101101 : data_out = 24'b000000000000001110000110;
    16'b1111011100101110 : data_out = 24'b000000000000001110000111;
    16'b1111011100101111 : data_out = 24'b000000000000001110000111;
    16'b1111011100110000 : data_out = 24'b000000000000001110001000;
    16'b1111011100110001 : data_out = 24'b000000000000001110001001;
    16'b1111011100110010 : data_out = 24'b000000000000001110001010;
    16'b1111011100110011 : data_out = 24'b000000000000001110001011;
    16'b1111011100110100 : data_out = 24'b000000000000001110001100;
    16'b1111011100110101 : data_out = 24'b000000000000001110001101;
    16'b1111011100110110 : data_out = 24'b000000000000001110001110;
    16'b1111011100110111 : data_out = 24'b000000000000001110001111;
    16'b1111011100111000 : data_out = 24'b000000000000001110001111;
    16'b1111011100111001 : data_out = 24'b000000000000001110010000;
    16'b1111011100111010 : data_out = 24'b000000000000001110010001;
    16'b1111011100111011 : data_out = 24'b000000000000001110010010;
    16'b1111011100111100 : data_out = 24'b000000000000001110010011;
    16'b1111011100111101 : data_out = 24'b000000000000001110010100;
    16'b1111011100111110 : data_out = 24'b000000000000001110010101;
    16'b1111011100111111 : data_out = 24'b000000000000001110010110;
    16'b1111011101000000 : data_out = 24'b000000000000001110010111;
    16'b1111011101000001 : data_out = 24'b000000000000001110011000;
    16'b1111011101000010 : data_out = 24'b000000000000001110011000;
    16'b1111011101000011 : data_out = 24'b000000000000001110011001;
    16'b1111011101000100 : data_out = 24'b000000000000001110011010;
    16'b1111011101000101 : data_out = 24'b000000000000001110011011;
    16'b1111011101000110 : data_out = 24'b000000000000001110011100;
    16'b1111011101000111 : data_out = 24'b000000000000001110011101;
    16'b1111011101001000 : data_out = 24'b000000000000001110011110;
    16'b1111011101001001 : data_out = 24'b000000000000001110011111;
    16'b1111011101001010 : data_out = 24'b000000000000001110100000;
    16'b1111011101001011 : data_out = 24'b000000000000001110100001;
    16'b1111011101001100 : data_out = 24'b000000000000001110100001;
    16'b1111011101001101 : data_out = 24'b000000000000001110100010;
    16'b1111011101001110 : data_out = 24'b000000000000001110100011;
    16'b1111011101001111 : data_out = 24'b000000000000001110100100;
    16'b1111011101010000 : data_out = 24'b000000000000001110100101;
    16'b1111011101010001 : data_out = 24'b000000000000001110100110;
    16'b1111011101010010 : data_out = 24'b000000000000001110100111;
    16'b1111011101010011 : data_out = 24'b000000000000001110101000;
    16'b1111011101010100 : data_out = 24'b000000000000001110101001;
    16'b1111011101010101 : data_out = 24'b000000000000001110101010;
    16'b1111011101010110 : data_out = 24'b000000000000001110101011;
    16'b1111011101010111 : data_out = 24'b000000000000001110101011;
    16'b1111011101011000 : data_out = 24'b000000000000001110101100;
    16'b1111011101011001 : data_out = 24'b000000000000001110101101;
    16'b1111011101011010 : data_out = 24'b000000000000001110101110;
    16'b1111011101011011 : data_out = 24'b000000000000001110101111;
    16'b1111011101011100 : data_out = 24'b000000000000001110110000;
    16'b1111011101011101 : data_out = 24'b000000000000001110110001;
    16'b1111011101011110 : data_out = 24'b000000000000001110110010;
    16'b1111011101011111 : data_out = 24'b000000000000001110110011;
    16'b1111011101100000 : data_out = 24'b000000000000001110110100;
    16'b1111011101100001 : data_out = 24'b000000000000001110110101;
    16'b1111011101100010 : data_out = 24'b000000000000001110110110;
    16'b1111011101100011 : data_out = 24'b000000000000001110110111;
    16'b1111011101100100 : data_out = 24'b000000000000001110111000;
    16'b1111011101100101 : data_out = 24'b000000000000001110111000;
    16'b1111011101100110 : data_out = 24'b000000000000001110111001;
    16'b1111011101100111 : data_out = 24'b000000000000001110111010;
    16'b1111011101101000 : data_out = 24'b000000000000001110111011;
    16'b1111011101101001 : data_out = 24'b000000000000001110111100;
    16'b1111011101101010 : data_out = 24'b000000000000001110111101;
    16'b1111011101101011 : data_out = 24'b000000000000001110111110;
    16'b1111011101101100 : data_out = 24'b000000000000001110111111;
    16'b1111011101101101 : data_out = 24'b000000000000001111000000;
    16'b1111011101101110 : data_out = 24'b000000000000001111000001;
    16'b1111011101101111 : data_out = 24'b000000000000001111000010;
    16'b1111011101110000 : data_out = 24'b000000000000001111000011;
    16'b1111011101110001 : data_out = 24'b000000000000001111000100;
    16'b1111011101110010 : data_out = 24'b000000000000001111000101;
    16'b1111011101110011 : data_out = 24'b000000000000001111000110;
    16'b1111011101110100 : data_out = 24'b000000000000001111000110;
    16'b1111011101110101 : data_out = 24'b000000000000001111000111;
    16'b1111011101110110 : data_out = 24'b000000000000001111001000;
    16'b1111011101110111 : data_out = 24'b000000000000001111001001;
    16'b1111011101111000 : data_out = 24'b000000000000001111001010;
    16'b1111011101111001 : data_out = 24'b000000000000001111001011;
    16'b1111011101111010 : data_out = 24'b000000000000001111001100;
    16'b1111011101111011 : data_out = 24'b000000000000001111001101;
    16'b1111011101111100 : data_out = 24'b000000000000001111001110;
    16'b1111011101111101 : data_out = 24'b000000000000001111001111;
    16'b1111011101111110 : data_out = 24'b000000000000001111010000;
    16'b1111011101111111 : data_out = 24'b000000000000001111010001;
    16'b1111011110000000 : data_out = 24'b000000000000001111010010;
    16'b1111011110000001 : data_out = 24'b000000000000001111010011;
    16'b1111011110000010 : data_out = 24'b000000000000001111010100;
    16'b1111011110000011 : data_out = 24'b000000000000001111010101;
    16'b1111011110000100 : data_out = 24'b000000000000001111010110;
    16'b1111011110000101 : data_out = 24'b000000000000001111010111;
    16'b1111011110000110 : data_out = 24'b000000000000001111011000;
    16'b1111011110000111 : data_out = 24'b000000000000001111011001;
    16'b1111011110001000 : data_out = 24'b000000000000001111011010;
    16'b1111011110001001 : data_out = 24'b000000000000001111011011;
    16'b1111011110001010 : data_out = 24'b000000000000001111011011;
    16'b1111011110001011 : data_out = 24'b000000000000001111011100;
    16'b1111011110001100 : data_out = 24'b000000000000001111011101;
    16'b1111011110001101 : data_out = 24'b000000000000001111011110;
    16'b1111011110001110 : data_out = 24'b000000000000001111011111;
    16'b1111011110001111 : data_out = 24'b000000000000001111100000;
    16'b1111011110010000 : data_out = 24'b000000000000001111100001;
    16'b1111011110010001 : data_out = 24'b000000000000001111100010;
    16'b1111011110010010 : data_out = 24'b000000000000001111100011;
    16'b1111011110010011 : data_out = 24'b000000000000001111100100;
    16'b1111011110010100 : data_out = 24'b000000000000001111100101;
    16'b1111011110010101 : data_out = 24'b000000000000001111100110;
    16'b1111011110010110 : data_out = 24'b000000000000001111100111;
    16'b1111011110010111 : data_out = 24'b000000000000001111101000;
    16'b1111011110011000 : data_out = 24'b000000000000001111101001;
    16'b1111011110011001 : data_out = 24'b000000000000001111101010;
    16'b1111011110011010 : data_out = 24'b000000000000001111101011;
    16'b1111011110011011 : data_out = 24'b000000000000001111101100;
    16'b1111011110011100 : data_out = 24'b000000000000001111101101;
    16'b1111011110011101 : data_out = 24'b000000000000001111101110;
    16'b1111011110011110 : data_out = 24'b000000000000001111101111;
    16'b1111011110011111 : data_out = 24'b000000000000001111110000;
    16'b1111011110100000 : data_out = 24'b000000000000001111110001;
    16'b1111011110100001 : data_out = 24'b000000000000001111110010;
    16'b1111011110100010 : data_out = 24'b000000000000001111110011;
    16'b1111011110100011 : data_out = 24'b000000000000001111110100;
    16'b1111011110100100 : data_out = 24'b000000000000001111110101;
    16'b1111011110100101 : data_out = 24'b000000000000001111110110;
    16'b1111011110100110 : data_out = 24'b000000000000001111110111;
    16'b1111011110100111 : data_out = 24'b000000000000001111111000;
    16'b1111011110101000 : data_out = 24'b000000000000001111111001;
    16'b1111011110101001 : data_out = 24'b000000000000001111111010;
    16'b1111011110101010 : data_out = 24'b000000000000001111111011;
    16'b1111011110101011 : data_out = 24'b000000000000001111111100;
    16'b1111011110101100 : data_out = 24'b000000000000001111111101;
    16'b1111011110101101 : data_out = 24'b000000000000001111111110;
    16'b1111011110101110 : data_out = 24'b000000000000001111111111;
    16'b1111011110101111 : data_out = 24'b000000000000010000000000;
    16'b1111011110110000 : data_out = 24'b000000000000010000000001;
    16'b1111011110110001 : data_out = 24'b000000000000010000000010;
    16'b1111011110110010 : data_out = 24'b000000000000010000000011;
    16'b1111011110110011 : data_out = 24'b000000000000010000000100;
    16'b1111011110110100 : data_out = 24'b000000000000010000000101;
    16'b1111011110110101 : data_out = 24'b000000000000010000000110;
    16'b1111011110110110 : data_out = 24'b000000000000010000000111;
    16'b1111011110110111 : data_out = 24'b000000000000010000001000;
    16'b1111011110111000 : data_out = 24'b000000000000010000001001;
    16'b1111011110111001 : data_out = 24'b000000000000010000001010;
    16'b1111011110111010 : data_out = 24'b000000000000010000001011;
    16'b1111011110111011 : data_out = 24'b000000000000010000001100;
    16'b1111011110111100 : data_out = 24'b000000000000010000001101;
    16'b1111011110111101 : data_out = 24'b000000000000010000001110;
    16'b1111011110111110 : data_out = 24'b000000000000010000001111;
    16'b1111011110111111 : data_out = 24'b000000000000010000010000;
    16'b1111011111000000 : data_out = 24'b000000000000010000010001;
    16'b1111011111000001 : data_out = 24'b000000000000010000010010;
    16'b1111011111000010 : data_out = 24'b000000000000010000010011;
    16'b1111011111000011 : data_out = 24'b000000000000010000010100;
    16'b1111011111000100 : data_out = 24'b000000000000010000010101;
    16'b1111011111000101 : data_out = 24'b000000000000010000010110;
    16'b1111011111000110 : data_out = 24'b000000000000010000010111;
    16'b1111011111000111 : data_out = 24'b000000000000010000011000;
    16'b1111011111001000 : data_out = 24'b000000000000010000011001;
    16'b1111011111001001 : data_out = 24'b000000000000010000011010;
    16'b1111011111001010 : data_out = 24'b000000000000010000011011;
    16'b1111011111001011 : data_out = 24'b000000000000010000011100;
    16'b1111011111001100 : data_out = 24'b000000000000010000011101;
    16'b1111011111001101 : data_out = 24'b000000000000010000011110;
    16'b1111011111001110 : data_out = 24'b000000000000010000011111;
    16'b1111011111001111 : data_out = 24'b000000000000010000100000;
    16'b1111011111010000 : data_out = 24'b000000000000010000100001;
    16'b1111011111010001 : data_out = 24'b000000000000010000100010;
    16'b1111011111010010 : data_out = 24'b000000000000010000100011;
    16'b1111011111010011 : data_out = 24'b000000000000010000100101;
    16'b1111011111010100 : data_out = 24'b000000000000010000100110;
    16'b1111011111010101 : data_out = 24'b000000000000010000100111;
    16'b1111011111010110 : data_out = 24'b000000000000010000101000;
    16'b1111011111010111 : data_out = 24'b000000000000010000101001;
    16'b1111011111011000 : data_out = 24'b000000000000010000101010;
    16'b1111011111011001 : data_out = 24'b000000000000010000101011;
    16'b1111011111011010 : data_out = 24'b000000000000010000101100;
    16'b1111011111011011 : data_out = 24'b000000000000010000101101;
    16'b1111011111011100 : data_out = 24'b000000000000010000101110;
    16'b1111011111011101 : data_out = 24'b000000000000010000101111;
    16'b1111011111011110 : data_out = 24'b000000000000010000110000;
    16'b1111011111011111 : data_out = 24'b000000000000010000110001;
    16'b1111011111100000 : data_out = 24'b000000000000010000110010;
    16'b1111011111100001 : data_out = 24'b000000000000010000110011;
    16'b1111011111100010 : data_out = 24'b000000000000010000110100;
    16'b1111011111100011 : data_out = 24'b000000000000010000110101;
    16'b1111011111100100 : data_out = 24'b000000000000010000110110;
    16'b1111011111100101 : data_out = 24'b000000000000010000110111;
    16'b1111011111100110 : data_out = 24'b000000000000010000111000;
    16'b1111011111100111 : data_out = 24'b000000000000010000111001;
    16'b1111011111101000 : data_out = 24'b000000000000010000111010;
    16'b1111011111101001 : data_out = 24'b000000000000010000111100;
    16'b1111011111101010 : data_out = 24'b000000000000010000111101;
    16'b1111011111101011 : data_out = 24'b000000000000010000111110;
    16'b1111011111101100 : data_out = 24'b000000000000010000111111;
    16'b1111011111101101 : data_out = 24'b000000000000010001000000;
    16'b1111011111101110 : data_out = 24'b000000000000010001000001;
    16'b1111011111101111 : data_out = 24'b000000000000010001000010;
    16'b1111011111110000 : data_out = 24'b000000000000010001000011;
    16'b1111011111110001 : data_out = 24'b000000000000010001000100;
    16'b1111011111110010 : data_out = 24'b000000000000010001000101;
    16'b1111011111110011 : data_out = 24'b000000000000010001000110;
    16'b1111011111110100 : data_out = 24'b000000000000010001000111;
    16'b1111011111110101 : data_out = 24'b000000000000010001001000;
    16'b1111011111110110 : data_out = 24'b000000000000010001001001;
    16'b1111011111110111 : data_out = 24'b000000000000010001001010;
    16'b1111011111111000 : data_out = 24'b000000000000010001001100;
    16'b1111011111111001 : data_out = 24'b000000000000010001001101;
    16'b1111011111111010 : data_out = 24'b000000000000010001001110;
    16'b1111011111111011 : data_out = 24'b000000000000010001001111;
    16'b1111011111111100 : data_out = 24'b000000000000010001010000;
    16'b1111011111111101 : data_out = 24'b000000000000010001010001;
    16'b1111011111111110 : data_out = 24'b000000000000010001010010;
    16'b1111011111111111 : data_out = 24'b000000000000010001010011;
    16'b1111100000000000 : data_out = 24'b000000000000010001010100;
    16'b1111100000000001 : data_out = 24'b000000000000010001010101;
    16'b1111100000000010 : data_out = 24'b000000000000010001010110;
    16'b1111100000000011 : data_out = 24'b000000000000010001010111;
    16'b1111100000000100 : data_out = 24'b000000000000010001011001;
    16'b1111100000000101 : data_out = 24'b000000000000010001011010;
    16'b1111100000000110 : data_out = 24'b000000000000010001011011;
    16'b1111100000000111 : data_out = 24'b000000000000010001011100;
    16'b1111100000001000 : data_out = 24'b000000000000010001011101;
    16'b1111100000001001 : data_out = 24'b000000000000010001011110;
    16'b1111100000001010 : data_out = 24'b000000000000010001011111;
    16'b1111100000001011 : data_out = 24'b000000000000010001100000;
    16'b1111100000001100 : data_out = 24'b000000000000010001100001;
    16'b1111100000001101 : data_out = 24'b000000000000010001100010;
    16'b1111100000001110 : data_out = 24'b000000000000010001100011;
    16'b1111100000001111 : data_out = 24'b000000000000010001100101;
    16'b1111100000010000 : data_out = 24'b000000000000010001100110;
    16'b1111100000010001 : data_out = 24'b000000000000010001100111;
    16'b1111100000010010 : data_out = 24'b000000000000010001101000;
    16'b1111100000010011 : data_out = 24'b000000000000010001101001;
    16'b1111100000010100 : data_out = 24'b000000000000010001101010;
    16'b1111100000010101 : data_out = 24'b000000000000010001101011;
    16'b1111100000010110 : data_out = 24'b000000000000010001101100;
    16'b1111100000010111 : data_out = 24'b000000000000010001101101;
    16'b1111100000011000 : data_out = 24'b000000000000010001101110;
    16'b1111100000011001 : data_out = 24'b000000000000010001110000;
    16'b1111100000011010 : data_out = 24'b000000000000010001110001;
    16'b1111100000011011 : data_out = 24'b000000000000010001110010;
    16'b1111100000011100 : data_out = 24'b000000000000010001110011;
    16'b1111100000011101 : data_out = 24'b000000000000010001110100;
    16'b1111100000011110 : data_out = 24'b000000000000010001110101;
    16'b1111100000011111 : data_out = 24'b000000000000010001110110;
    16'b1111100000100000 : data_out = 24'b000000000000010001110111;
    16'b1111100000100001 : data_out = 24'b000000000000010001111000;
    16'b1111100000100010 : data_out = 24'b000000000000010001111010;
    16'b1111100000100011 : data_out = 24'b000000000000010001111011;
    16'b1111100000100100 : data_out = 24'b000000000000010001111100;
    16'b1111100000100101 : data_out = 24'b000000000000010001111101;
    16'b1111100000100110 : data_out = 24'b000000000000010001111110;
    16'b1111100000100111 : data_out = 24'b000000000000010001111111;
    16'b1111100000101000 : data_out = 24'b000000000000010010000000;
    16'b1111100000101001 : data_out = 24'b000000000000010010000001;
    16'b1111100000101010 : data_out = 24'b000000000000010010000011;
    16'b1111100000101011 : data_out = 24'b000000000000010010000100;
    16'b1111100000101100 : data_out = 24'b000000000000010010000101;
    16'b1111100000101101 : data_out = 24'b000000000000010010000110;
    16'b1111100000101110 : data_out = 24'b000000000000010010000111;
    16'b1111100000101111 : data_out = 24'b000000000000010010001000;
    16'b1111100000110000 : data_out = 24'b000000000000010010001001;
    16'b1111100000110001 : data_out = 24'b000000000000010010001011;
    16'b1111100000110010 : data_out = 24'b000000000000010010001100;
    16'b1111100000110011 : data_out = 24'b000000000000010010001101;
    16'b1111100000110100 : data_out = 24'b000000000000010010001110;
    16'b1111100000110101 : data_out = 24'b000000000000010010001111;
    16'b1111100000110110 : data_out = 24'b000000000000010010010000;
    16'b1111100000110111 : data_out = 24'b000000000000010010010001;
    16'b1111100000111000 : data_out = 24'b000000000000010010010010;
    16'b1111100000111001 : data_out = 24'b000000000000010010010100;
    16'b1111100000111010 : data_out = 24'b000000000000010010010101;
    16'b1111100000111011 : data_out = 24'b000000000000010010010110;
    16'b1111100000111100 : data_out = 24'b000000000000010010010111;
    16'b1111100000111101 : data_out = 24'b000000000000010010011000;
    16'b1111100000111110 : data_out = 24'b000000000000010010011001;
    16'b1111100000111111 : data_out = 24'b000000000000010010011011;
    16'b1111100001000000 : data_out = 24'b000000000000010010011100;
    16'b1111100001000001 : data_out = 24'b000000000000010010011101;
    16'b1111100001000010 : data_out = 24'b000000000000010010011110;
    16'b1111100001000011 : data_out = 24'b000000000000010010011111;
    16'b1111100001000100 : data_out = 24'b000000000000010010100000;
    16'b1111100001000101 : data_out = 24'b000000000000010010100001;
    16'b1111100001000110 : data_out = 24'b000000000000010010100011;
    16'b1111100001000111 : data_out = 24'b000000000000010010100100;
    16'b1111100001001000 : data_out = 24'b000000000000010010100101;
    16'b1111100001001001 : data_out = 24'b000000000000010010100110;
    16'b1111100001001010 : data_out = 24'b000000000000010010100111;
    16'b1111100001001011 : data_out = 24'b000000000000010010101000;
    16'b1111100001001100 : data_out = 24'b000000000000010010101010;
    16'b1111100001001101 : data_out = 24'b000000000000010010101011;
    16'b1111100001001110 : data_out = 24'b000000000000010010101100;
    16'b1111100001001111 : data_out = 24'b000000000000010010101101;
    16'b1111100001010000 : data_out = 24'b000000000000010010101110;
    16'b1111100001010001 : data_out = 24'b000000000000010010101111;
    16'b1111100001010010 : data_out = 24'b000000000000010010110001;
    16'b1111100001010011 : data_out = 24'b000000000000010010110010;
    16'b1111100001010100 : data_out = 24'b000000000000010010110011;
    16'b1111100001010101 : data_out = 24'b000000000000010010110100;
    16'b1111100001010110 : data_out = 24'b000000000000010010110101;
    16'b1111100001010111 : data_out = 24'b000000000000010010110110;
    16'b1111100001011000 : data_out = 24'b000000000000010010111000;
    16'b1111100001011001 : data_out = 24'b000000000000010010111001;
    16'b1111100001011010 : data_out = 24'b000000000000010010111010;
    16'b1111100001011011 : data_out = 24'b000000000000010010111011;
    16'b1111100001011100 : data_out = 24'b000000000000010010111100;
    16'b1111100001011101 : data_out = 24'b000000000000010010111110;
    16'b1111100001011110 : data_out = 24'b000000000000010010111111;
    16'b1111100001011111 : data_out = 24'b000000000000010011000000;
    16'b1111100001100000 : data_out = 24'b000000000000010011000001;
    16'b1111100001100001 : data_out = 24'b000000000000010011000010;
    16'b1111100001100010 : data_out = 24'b000000000000010011000100;
    16'b1111100001100011 : data_out = 24'b000000000000010011000101;
    16'b1111100001100100 : data_out = 24'b000000000000010011000110;
    16'b1111100001100101 : data_out = 24'b000000000000010011000111;
    16'b1111100001100110 : data_out = 24'b000000000000010011001000;
    16'b1111100001100111 : data_out = 24'b000000000000010011001001;
    16'b1111100001101000 : data_out = 24'b000000000000010011001011;
    16'b1111100001101001 : data_out = 24'b000000000000010011001100;
    16'b1111100001101010 : data_out = 24'b000000000000010011001101;
    16'b1111100001101011 : data_out = 24'b000000000000010011001110;
    16'b1111100001101100 : data_out = 24'b000000000000010011001111;
    16'b1111100001101101 : data_out = 24'b000000000000010011010001;
    16'b1111100001101110 : data_out = 24'b000000000000010011010010;
    16'b1111100001101111 : data_out = 24'b000000000000010011010011;
    16'b1111100001110000 : data_out = 24'b000000000000010011010100;
    16'b1111100001110001 : data_out = 24'b000000000000010011010110;
    16'b1111100001110010 : data_out = 24'b000000000000010011010111;
    16'b1111100001110011 : data_out = 24'b000000000000010011011000;
    16'b1111100001110100 : data_out = 24'b000000000000010011011001;
    16'b1111100001110101 : data_out = 24'b000000000000010011011010;
    16'b1111100001110110 : data_out = 24'b000000000000010011011100;
    16'b1111100001110111 : data_out = 24'b000000000000010011011101;
    16'b1111100001111000 : data_out = 24'b000000000000010011011110;
    16'b1111100001111001 : data_out = 24'b000000000000010011011111;
    16'b1111100001111010 : data_out = 24'b000000000000010011100000;
    16'b1111100001111011 : data_out = 24'b000000000000010011100010;
    16'b1111100001111100 : data_out = 24'b000000000000010011100011;
    16'b1111100001111101 : data_out = 24'b000000000000010011100100;
    16'b1111100001111110 : data_out = 24'b000000000000010011100101;
    16'b1111100001111111 : data_out = 24'b000000000000010011100111;
    16'b1111100010000000 : data_out = 24'b000000000000010011101000;
    16'b1111100010000001 : data_out = 24'b000000000000010011101001;
    16'b1111100010000010 : data_out = 24'b000000000000010011101010;
    16'b1111100010000011 : data_out = 24'b000000000000010011101011;
    16'b1111100010000100 : data_out = 24'b000000000000010011101101;
    16'b1111100010000101 : data_out = 24'b000000000000010011101110;
    16'b1111100010000110 : data_out = 24'b000000000000010011101111;
    16'b1111100010000111 : data_out = 24'b000000000000010011110000;
    16'b1111100010001000 : data_out = 24'b000000000000010011110010;
    16'b1111100010001001 : data_out = 24'b000000000000010011110011;
    16'b1111100010001010 : data_out = 24'b000000000000010011110100;
    16'b1111100010001011 : data_out = 24'b000000000000010011110101;
    16'b1111100010001100 : data_out = 24'b000000000000010011110111;
    16'b1111100010001101 : data_out = 24'b000000000000010011111000;
    16'b1111100010001110 : data_out = 24'b000000000000010011111001;
    16'b1111100010001111 : data_out = 24'b000000000000010011111010;
    16'b1111100010010000 : data_out = 24'b000000000000010011111100;
    16'b1111100010010001 : data_out = 24'b000000000000010011111101;
    16'b1111100010010010 : data_out = 24'b000000000000010011111110;
    16'b1111100010010011 : data_out = 24'b000000000000010011111111;
    16'b1111100010010100 : data_out = 24'b000000000000010100000001;
    16'b1111100010010101 : data_out = 24'b000000000000010100000010;
    16'b1111100010010110 : data_out = 24'b000000000000010100000011;
    16'b1111100010010111 : data_out = 24'b000000000000010100000100;
    16'b1111100010011000 : data_out = 24'b000000000000010100000110;
    16'b1111100010011001 : data_out = 24'b000000000000010100000111;
    16'b1111100010011010 : data_out = 24'b000000000000010100001000;
    16'b1111100010011011 : data_out = 24'b000000000000010100001001;
    16'b1111100010011100 : data_out = 24'b000000000000010100001011;
    16'b1111100010011101 : data_out = 24'b000000000000010100001100;
    16'b1111100010011110 : data_out = 24'b000000000000010100001101;
    16'b1111100010011111 : data_out = 24'b000000000000010100001110;
    16'b1111100010100000 : data_out = 24'b000000000000010100010000;
    16'b1111100010100001 : data_out = 24'b000000000000010100010001;
    16'b1111100010100010 : data_out = 24'b000000000000010100010010;
    16'b1111100010100011 : data_out = 24'b000000000000010100010011;
    16'b1111100010100100 : data_out = 24'b000000000000010100010101;
    16'b1111100010100101 : data_out = 24'b000000000000010100010110;
    16'b1111100010100110 : data_out = 24'b000000000000010100010111;
    16'b1111100010100111 : data_out = 24'b000000000000010100011001;
    16'b1111100010101000 : data_out = 24'b000000000000010100011010;
    16'b1111100010101001 : data_out = 24'b000000000000010100011011;
    16'b1111100010101010 : data_out = 24'b000000000000010100011100;
    16'b1111100010101011 : data_out = 24'b000000000000010100011110;
    16'b1111100010101100 : data_out = 24'b000000000000010100011111;
    16'b1111100010101101 : data_out = 24'b000000000000010100100000;
    16'b1111100010101110 : data_out = 24'b000000000000010100100010;
    16'b1111100010101111 : data_out = 24'b000000000000010100100011;
    16'b1111100010110000 : data_out = 24'b000000000000010100100100;
    16'b1111100010110001 : data_out = 24'b000000000000010100100101;
    16'b1111100010110010 : data_out = 24'b000000000000010100100111;
    16'b1111100010110011 : data_out = 24'b000000000000010100101000;
    16'b1111100010110100 : data_out = 24'b000000000000010100101001;
    16'b1111100010110101 : data_out = 24'b000000000000010100101011;
    16'b1111100010110110 : data_out = 24'b000000000000010100101100;
    16'b1111100010110111 : data_out = 24'b000000000000010100101101;
    16'b1111100010111000 : data_out = 24'b000000000000010100101110;
    16'b1111100010111001 : data_out = 24'b000000000000010100110000;
    16'b1111100010111010 : data_out = 24'b000000000000010100110001;
    16'b1111100010111011 : data_out = 24'b000000000000010100110010;
    16'b1111100010111100 : data_out = 24'b000000000000010100110100;
    16'b1111100010111101 : data_out = 24'b000000000000010100110101;
    16'b1111100010111110 : data_out = 24'b000000000000010100110110;
    16'b1111100010111111 : data_out = 24'b000000000000010100111000;
    16'b1111100011000000 : data_out = 24'b000000000000010100111001;
    16'b1111100011000001 : data_out = 24'b000000000000010100111010;
    16'b1111100011000010 : data_out = 24'b000000000000010100111011;
    16'b1111100011000011 : data_out = 24'b000000000000010100111101;
    16'b1111100011000100 : data_out = 24'b000000000000010100111110;
    16'b1111100011000101 : data_out = 24'b000000000000010100111111;
    16'b1111100011000110 : data_out = 24'b000000000000010101000001;
    16'b1111100011000111 : data_out = 24'b000000000000010101000010;
    16'b1111100011001000 : data_out = 24'b000000000000010101000011;
    16'b1111100011001001 : data_out = 24'b000000000000010101000101;
    16'b1111100011001010 : data_out = 24'b000000000000010101000110;
    16'b1111100011001011 : data_out = 24'b000000000000010101000111;
    16'b1111100011001100 : data_out = 24'b000000000000010101001001;
    16'b1111100011001101 : data_out = 24'b000000000000010101001010;
    16'b1111100011001110 : data_out = 24'b000000000000010101001011;
    16'b1111100011001111 : data_out = 24'b000000000000010101001101;
    16'b1111100011010000 : data_out = 24'b000000000000010101001110;
    16'b1111100011010001 : data_out = 24'b000000000000010101001111;
    16'b1111100011010010 : data_out = 24'b000000000000010101010001;
    16'b1111100011010011 : data_out = 24'b000000000000010101010010;
    16'b1111100011010100 : data_out = 24'b000000000000010101010011;
    16'b1111100011010101 : data_out = 24'b000000000000010101010101;
    16'b1111100011010110 : data_out = 24'b000000000000010101010110;
    16'b1111100011010111 : data_out = 24'b000000000000010101010111;
    16'b1111100011011000 : data_out = 24'b000000000000010101011001;
    16'b1111100011011001 : data_out = 24'b000000000000010101011010;
    16'b1111100011011010 : data_out = 24'b000000000000010101011011;
    16'b1111100011011011 : data_out = 24'b000000000000010101011101;
    16'b1111100011011100 : data_out = 24'b000000000000010101011110;
    16'b1111100011011101 : data_out = 24'b000000000000010101011111;
    16'b1111100011011110 : data_out = 24'b000000000000010101100001;
    16'b1111100011011111 : data_out = 24'b000000000000010101100010;
    16'b1111100011100000 : data_out = 24'b000000000000010101100011;
    16'b1111100011100001 : data_out = 24'b000000000000010101100101;
    16'b1111100011100010 : data_out = 24'b000000000000010101100110;
    16'b1111100011100011 : data_out = 24'b000000000000010101100111;
    16'b1111100011100100 : data_out = 24'b000000000000010101101001;
    16'b1111100011100101 : data_out = 24'b000000000000010101101010;
    16'b1111100011100110 : data_out = 24'b000000000000010101101011;
    16'b1111100011100111 : data_out = 24'b000000000000010101101101;
    16'b1111100011101000 : data_out = 24'b000000000000010101101110;
    16'b1111100011101001 : data_out = 24'b000000000000010101101111;
    16'b1111100011101010 : data_out = 24'b000000000000010101110001;
    16'b1111100011101011 : data_out = 24'b000000000000010101110010;
    16'b1111100011101100 : data_out = 24'b000000000000010101110100;
    16'b1111100011101101 : data_out = 24'b000000000000010101110101;
    16'b1111100011101110 : data_out = 24'b000000000000010101110110;
    16'b1111100011101111 : data_out = 24'b000000000000010101111000;
    16'b1111100011110000 : data_out = 24'b000000000000010101111001;
    16'b1111100011110001 : data_out = 24'b000000000000010101111010;
    16'b1111100011110010 : data_out = 24'b000000000000010101111100;
    16'b1111100011110011 : data_out = 24'b000000000000010101111101;
    16'b1111100011110100 : data_out = 24'b000000000000010101111110;
    16'b1111100011110101 : data_out = 24'b000000000000010110000000;
    16'b1111100011110110 : data_out = 24'b000000000000010110000001;
    16'b1111100011110111 : data_out = 24'b000000000000010110000011;
    16'b1111100011111000 : data_out = 24'b000000000000010110000100;
    16'b1111100011111001 : data_out = 24'b000000000000010110000101;
    16'b1111100011111010 : data_out = 24'b000000000000010110000111;
    16'b1111100011111011 : data_out = 24'b000000000000010110001000;
    16'b1111100011111100 : data_out = 24'b000000000000010110001010;
    16'b1111100011111101 : data_out = 24'b000000000000010110001011;
    16'b1111100011111110 : data_out = 24'b000000000000010110001100;
    16'b1111100011111111 : data_out = 24'b000000000000010110001110;
    16'b1111100100000000 : data_out = 24'b000000000000010110001111;
    16'b1111100100000001 : data_out = 24'b000000000000010110010000;
    16'b1111100100000010 : data_out = 24'b000000000000010110010010;
    16'b1111100100000011 : data_out = 24'b000000000000010110010011;
    16'b1111100100000100 : data_out = 24'b000000000000010110010101;
    16'b1111100100000101 : data_out = 24'b000000000000010110010110;
    16'b1111100100000110 : data_out = 24'b000000000000010110010111;
    16'b1111100100000111 : data_out = 24'b000000000000010110011001;
    16'b1111100100001000 : data_out = 24'b000000000000010110011010;
    16'b1111100100001001 : data_out = 24'b000000000000010110011100;
    16'b1111100100001010 : data_out = 24'b000000000000010110011101;
    16'b1111100100001011 : data_out = 24'b000000000000010110011110;
    16'b1111100100001100 : data_out = 24'b000000000000010110100000;
    16'b1111100100001101 : data_out = 24'b000000000000010110100001;
    16'b1111100100001110 : data_out = 24'b000000000000010110100011;
    16'b1111100100001111 : data_out = 24'b000000000000010110100100;
    16'b1111100100010000 : data_out = 24'b000000000000010110100101;
    16'b1111100100010001 : data_out = 24'b000000000000010110100111;
    16'b1111100100010010 : data_out = 24'b000000000000010110101000;
    16'b1111100100010011 : data_out = 24'b000000000000010110101010;
    16'b1111100100010100 : data_out = 24'b000000000000010110101011;
    16'b1111100100010101 : data_out = 24'b000000000000010110101101;
    16'b1111100100010110 : data_out = 24'b000000000000010110101110;
    16'b1111100100010111 : data_out = 24'b000000000000010110101111;
    16'b1111100100011000 : data_out = 24'b000000000000010110110001;
    16'b1111100100011001 : data_out = 24'b000000000000010110110010;
    16'b1111100100011010 : data_out = 24'b000000000000010110110100;
    16'b1111100100011011 : data_out = 24'b000000000000010110110101;
    16'b1111100100011100 : data_out = 24'b000000000000010110110111;
    16'b1111100100011101 : data_out = 24'b000000000000010110111000;
    16'b1111100100011110 : data_out = 24'b000000000000010110111001;
    16'b1111100100011111 : data_out = 24'b000000000000010110111011;
    16'b1111100100100000 : data_out = 24'b000000000000010110111100;
    16'b1111100100100001 : data_out = 24'b000000000000010110111110;
    16'b1111100100100010 : data_out = 24'b000000000000010110111111;
    16'b1111100100100011 : data_out = 24'b000000000000010111000001;
    16'b1111100100100100 : data_out = 24'b000000000000010111000010;
    16'b1111100100100101 : data_out = 24'b000000000000010111000011;
    16'b1111100100100110 : data_out = 24'b000000000000010111000101;
    16'b1111100100100111 : data_out = 24'b000000000000010111000110;
    16'b1111100100101000 : data_out = 24'b000000000000010111001000;
    16'b1111100100101001 : data_out = 24'b000000000000010111001001;
    16'b1111100100101010 : data_out = 24'b000000000000010111001011;
    16'b1111100100101011 : data_out = 24'b000000000000010111001100;
    16'b1111100100101100 : data_out = 24'b000000000000010111001110;
    16'b1111100100101101 : data_out = 24'b000000000000010111001111;
    16'b1111100100101110 : data_out = 24'b000000000000010111010000;
    16'b1111100100101111 : data_out = 24'b000000000000010111010010;
    16'b1111100100110000 : data_out = 24'b000000000000010111010011;
    16'b1111100100110001 : data_out = 24'b000000000000010111010101;
    16'b1111100100110010 : data_out = 24'b000000000000010111010110;
    16'b1111100100110011 : data_out = 24'b000000000000010111011000;
    16'b1111100100110100 : data_out = 24'b000000000000010111011001;
    16'b1111100100110101 : data_out = 24'b000000000000010111011011;
    16'b1111100100110110 : data_out = 24'b000000000000010111011100;
    16'b1111100100110111 : data_out = 24'b000000000000010111011110;
    16'b1111100100111000 : data_out = 24'b000000000000010111011111;
    16'b1111100100111001 : data_out = 24'b000000000000010111100001;
    16'b1111100100111010 : data_out = 24'b000000000000010111100010;
    16'b1111100100111011 : data_out = 24'b000000000000010111100011;
    16'b1111100100111100 : data_out = 24'b000000000000010111100101;
    16'b1111100100111101 : data_out = 24'b000000000000010111100110;
    16'b1111100100111110 : data_out = 24'b000000000000010111101000;
    16'b1111100100111111 : data_out = 24'b000000000000010111101001;
    16'b1111100101000000 : data_out = 24'b000000000000010111101011;
    16'b1111100101000001 : data_out = 24'b000000000000010111101100;
    16'b1111100101000010 : data_out = 24'b000000000000010111101110;
    16'b1111100101000011 : data_out = 24'b000000000000010111101111;
    16'b1111100101000100 : data_out = 24'b000000000000010111110001;
    16'b1111100101000101 : data_out = 24'b000000000000010111110010;
    16'b1111100101000110 : data_out = 24'b000000000000010111110100;
    16'b1111100101000111 : data_out = 24'b000000000000010111110101;
    16'b1111100101001000 : data_out = 24'b000000000000010111110111;
    16'b1111100101001001 : data_out = 24'b000000000000010111111000;
    16'b1111100101001010 : data_out = 24'b000000000000010111111010;
    16'b1111100101001011 : data_out = 24'b000000000000010111111011;
    16'b1111100101001100 : data_out = 24'b000000000000010111111101;
    16'b1111100101001101 : data_out = 24'b000000000000010111111110;
    16'b1111100101001110 : data_out = 24'b000000000000011000000000;
    16'b1111100101001111 : data_out = 24'b000000000000011000000001;
    16'b1111100101010000 : data_out = 24'b000000000000011000000011;
    16'b1111100101010001 : data_out = 24'b000000000000011000000100;
    16'b1111100101010010 : data_out = 24'b000000000000011000000110;
    16'b1111100101010011 : data_out = 24'b000000000000011000000111;
    16'b1111100101010100 : data_out = 24'b000000000000011000001001;
    16'b1111100101010101 : data_out = 24'b000000000000011000001010;
    16'b1111100101010110 : data_out = 24'b000000000000011000001100;
    16'b1111100101010111 : data_out = 24'b000000000000011000001101;
    16'b1111100101011000 : data_out = 24'b000000000000011000001111;
    16'b1111100101011001 : data_out = 24'b000000000000011000010000;
    16'b1111100101011010 : data_out = 24'b000000000000011000010010;
    16'b1111100101011011 : data_out = 24'b000000000000011000010011;
    16'b1111100101011100 : data_out = 24'b000000000000011000010101;
    16'b1111100101011101 : data_out = 24'b000000000000011000010110;
    16'b1111100101011110 : data_out = 24'b000000000000011000011000;
    16'b1111100101011111 : data_out = 24'b000000000000011000011001;
    16'b1111100101100000 : data_out = 24'b000000000000011000011011;
    16'b1111100101100001 : data_out = 24'b000000000000011000011100;
    16'b1111100101100010 : data_out = 24'b000000000000011000011110;
    16'b1111100101100011 : data_out = 24'b000000000000011000100000;
    16'b1111100101100100 : data_out = 24'b000000000000011000100001;
    16'b1111100101100101 : data_out = 24'b000000000000011000100011;
    16'b1111100101100110 : data_out = 24'b000000000000011000100100;
    16'b1111100101100111 : data_out = 24'b000000000000011000100110;
    16'b1111100101101000 : data_out = 24'b000000000000011000100111;
    16'b1111100101101001 : data_out = 24'b000000000000011000101001;
    16'b1111100101101010 : data_out = 24'b000000000000011000101010;
    16'b1111100101101011 : data_out = 24'b000000000000011000101100;
    16'b1111100101101100 : data_out = 24'b000000000000011000101101;
    16'b1111100101101101 : data_out = 24'b000000000000011000101111;
    16'b1111100101101110 : data_out = 24'b000000000000011000110000;
    16'b1111100101101111 : data_out = 24'b000000000000011000110010;
    16'b1111100101110000 : data_out = 24'b000000000000011000110100;
    16'b1111100101110001 : data_out = 24'b000000000000011000110101;
    16'b1111100101110010 : data_out = 24'b000000000000011000110111;
    16'b1111100101110011 : data_out = 24'b000000000000011000111000;
    16'b1111100101110100 : data_out = 24'b000000000000011000111010;
    16'b1111100101110101 : data_out = 24'b000000000000011000111011;
    16'b1111100101110110 : data_out = 24'b000000000000011000111101;
    16'b1111100101110111 : data_out = 24'b000000000000011000111110;
    16'b1111100101111000 : data_out = 24'b000000000000011001000000;
    16'b1111100101111001 : data_out = 24'b000000000000011001000010;
    16'b1111100101111010 : data_out = 24'b000000000000011001000011;
    16'b1111100101111011 : data_out = 24'b000000000000011001000101;
    16'b1111100101111100 : data_out = 24'b000000000000011001000110;
    16'b1111100101111101 : data_out = 24'b000000000000011001001000;
    16'b1111100101111110 : data_out = 24'b000000000000011001001001;
    16'b1111100101111111 : data_out = 24'b000000000000011001001011;
    16'b1111100110000000 : data_out = 24'b000000000000011001001101;
    16'b1111100110000001 : data_out = 24'b000000000000011001001110;
    16'b1111100110000010 : data_out = 24'b000000000000011001010000;
    16'b1111100110000011 : data_out = 24'b000000000000011001010001;
    16'b1111100110000100 : data_out = 24'b000000000000011001010011;
    16'b1111100110000101 : data_out = 24'b000000000000011001010100;
    16'b1111100110000110 : data_out = 24'b000000000000011001010110;
    16'b1111100110000111 : data_out = 24'b000000000000011001011000;
    16'b1111100110001000 : data_out = 24'b000000000000011001011001;
    16'b1111100110001001 : data_out = 24'b000000000000011001011011;
    16'b1111100110001010 : data_out = 24'b000000000000011001011100;
    16'b1111100110001011 : data_out = 24'b000000000000011001011110;
    16'b1111100110001100 : data_out = 24'b000000000000011001100000;
    16'b1111100110001101 : data_out = 24'b000000000000011001100001;
    16'b1111100110001110 : data_out = 24'b000000000000011001100011;
    16'b1111100110001111 : data_out = 24'b000000000000011001100100;
    16'b1111100110010000 : data_out = 24'b000000000000011001100110;
    16'b1111100110010001 : data_out = 24'b000000000000011001101000;
    16'b1111100110010010 : data_out = 24'b000000000000011001101001;
    16'b1111100110010011 : data_out = 24'b000000000000011001101011;
    16'b1111100110010100 : data_out = 24'b000000000000011001101100;
    16'b1111100110010101 : data_out = 24'b000000000000011001101110;
    16'b1111100110010110 : data_out = 24'b000000000000011001110000;
    16'b1111100110010111 : data_out = 24'b000000000000011001110001;
    16'b1111100110011000 : data_out = 24'b000000000000011001110011;
    16'b1111100110011001 : data_out = 24'b000000000000011001110100;
    16'b1111100110011010 : data_out = 24'b000000000000011001110110;
    16'b1111100110011011 : data_out = 24'b000000000000011001111000;
    16'b1111100110011100 : data_out = 24'b000000000000011001111001;
    16'b1111100110011101 : data_out = 24'b000000000000011001111011;
    16'b1111100110011110 : data_out = 24'b000000000000011001111101;
    16'b1111100110011111 : data_out = 24'b000000000000011001111110;
    16'b1111100110100000 : data_out = 24'b000000000000011010000000;
    16'b1111100110100001 : data_out = 24'b000000000000011010000001;
    16'b1111100110100010 : data_out = 24'b000000000000011010000011;
    16'b1111100110100011 : data_out = 24'b000000000000011010000101;
    16'b1111100110100100 : data_out = 24'b000000000000011010000110;
    16'b1111100110100101 : data_out = 24'b000000000000011010001000;
    16'b1111100110100110 : data_out = 24'b000000000000011010001010;
    16'b1111100110100111 : data_out = 24'b000000000000011010001011;
    16'b1111100110101000 : data_out = 24'b000000000000011010001101;
    16'b1111100110101001 : data_out = 24'b000000000000011010001110;
    16'b1111100110101010 : data_out = 24'b000000000000011010010000;
    16'b1111100110101011 : data_out = 24'b000000000000011010010010;
    16'b1111100110101100 : data_out = 24'b000000000000011010010011;
    16'b1111100110101101 : data_out = 24'b000000000000011010010101;
    16'b1111100110101110 : data_out = 24'b000000000000011010010111;
    16'b1111100110101111 : data_out = 24'b000000000000011010011000;
    16'b1111100110110000 : data_out = 24'b000000000000011010011010;
    16'b1111100110110001 : data_out = 24'b000000000000011010011100;
    16'b1111100110110010 : data_out = 24'b000000000000011010011101;
    16'b1111100110110011 : data_out = 24'b000000000000011010011111;
    16'b1111100110110100 : data_out = 24'b000000000000011010100001;
    16'b1111100110110101 : data_out = 24'b000000000000011010100010;
    16'b1111100110110110 : data_out = 24'b000000000000011010100100;
    16'b1111100110110111 : data_out = 24'b000000000000011010100110;
    16'b1111100110111000 : data_out = 24'b000000000000011010100111;
    16'b1111100110111001 : data_out = 24'b000000000000011010101001;
    16'b1111100110111010 : data_out = 24'b000000000000011010101011;
    16'b1111100110111011 : data_out = 24'b000000000000011010101100;
    16'b1111100110111100 : data_out = 24'b000000000000011010101110;
    16'b1111100110111101 : data_out = 24'b000000000000011010110000;
    16'b1111100110111110 : data_out = 24'b000000000000011010110001;
    16'b1111100110111111 : data_out = 24'b000000000000011010110011;
    16'b1111100111000000 : data_out = 24'b000000000000011010110101;
    16'b1111100111000001 : data_out = 24'b000000000000011010110110;
    16'b1111100111000010 : data_out = 24'b000000000000011010111000;
    16'b1111100111000011 : data_out = 24'b000000000000011010111010;
    16'b1111100111000100 : data_out = 24'b000000000000011010111011;
    16'b1111100111000101 : data_out = 24'b000000000000011010111101;
    16'b1111100111000110 : data_out = 24'b000000000000011010111111;
    16'b1111100111000111 : data_out = 24'b000000000000011011000000;
    16'b1111100111001000 : data_out = 24'b000000000000011011000010;
    16'b1111100111001001 : data_out = 24'b000000000000011011000100;
    16'b1111100111001010 : data_out = 24'b000000000000011011000101;
    16'b1111100111001011 : data_out = 24'b000000000000011011000111;
    16'b1111100111001100 : data_out = 24'b000000000000011011001001;
    16'b1111100111001101 : data_out = 24'b000000000000011011001011;
    16'b1111100111001110 : data_out = 24'b000000000000011011001100;
    16'b1111100111001111 : data_out = 24'b000000000000011011001110;
    16'b1111100111010000 : data_out = 24'b000000000000011011010000;
    16'b1111100111010001 : data_out = 24'b000000000000011011010001;
    16'b1111100111010010 : data_out = 24'b000000000000011011010011;
    16'b1111100111010011 : data_out = 24'b000000000000011011010101;
    16'b1111100111010100 : data_out = 24'b000000000000011011010111;
    16'b1111100111010101 : data_out = 24'b000000000000011011011000;
    16'b1111100111010110 : data_out = 24'b000000000000011011011010;
    16'b1111100111010111 : data_out = 24'b000000000000011011011100;
    16'b1111100111011000 : data_out = 24'b000000000000011011011101;
    16'b1111100111011001 : data_out = 24'b000000000000011011011111;
    16'b1111100111011010 : data_out = 24'b000000000000011011100001;
    16'b1111100111011011 : data_out = 24'b000000000000011011100011;
    16'b1111100111011100 : data_out = 24'b000000000000011011100100;
    16'b1111100111011101 : data_out = 24'b000000000000011011100110;
    16'b1111100111011110 : data_out = 24'b000000000000011011101000;
    16'b1111100111011111 : data_out = 24'b000000000000011011101001;
    16'b1111100111100000 : data_out = 24'b000000000000011011101011;
    16'b1111100111100001 : data_out = 24'b000000000000011011101101;
    16'b1111100111100010 : data_out = 24'b000000000000011011101111;
    16'b1111100111100011 : data_out = 24'b000000000000011011110000;
    16'b1111100111100100 : data_out = 24'b000000000000011011110010;
    16'b1111100111100101 : data_out = 24'b000000000000011011110100;
    16'b1111100111100110 : data_out = 24'b000000000000011011110110;
    16'b1111100111100111 : data_out = 24'b000000000000011011110111;
    16'b1111100111101000 : data_out = 24'b000000000000011011111001;
    16'b1111100111101001 : data_out = 24'b000000000000011011111011;
    16'b1111100111101010 : data_out = 24'b000000000000011011111101;
    16'b1111100111101011 : data_out = 24'b000000000000011011111110;
    16'b1111100111101100 : data_out = 24'b000000000000011100000000;
    16'b1111100111101101 : data_out = 24'b000000000000011100000010;
    16'b1111100111101110 : data_out = 24'b000000000000011100000100;
    16'b1111100111101111 : data_out = 24'b000000000000011100000101;
    16'b1111100111110000 : data_out = 24'b000000000000011100000111;
    16'b1111100111110001 : data_out = 24'b000000000000011100001001;
    16'b1111100111110010 : data_out = 24'b000000000000011100001011;
    16'b1111100111110011 : data_out = 24'b000000000000011100001100;
    16'b1111100111110100 : data_out = 24'b000000000000011100001110;
    16'b1111100111110101 : data_out = 24'b000000000000011100010000;
    16'b1111100111110110 : data_out = 24'b000000000000011100010010;
    16'b1111100111110111 : data_out = 24'b000000000000011100010011;
    16'b1111100111111000 : data_out = 24'b000000000000011100010101;
    16'b1111100111111001 : data_out = 24'b000000000000011100010111;
    16'b1111100111111010 : data_out = 24'b000000000000011100011001;
    16'b1111100111111011 : data_out = 24'b000000000000011100011010;
    16'b1111100111111100 : data_out = 24'b000000000000011100011100;
    16'b1111100111111101 : data_out = 24'b000000000000011100011110;
    16'b1111100111111110 : data_out = 24'b000000000000011100100000;
    16'b1111100111111111 : data_out = 24'b000000000000011100100010;
    16'b1111101000000000 : data_out = 24'b000000000000011100100011;
    16'b1111101000000001 : data_out = 24'b000000000000011100100101;
    16'b1111101000000010 : data_out = 24'b000000000000011100100111;
    16'b1111101000000011 : data_out = 24'b000000000000011100101001;
    16'b1111101000000100 : data_out = 24'b000000000000011100101011;
    16'b1111101000000101 : data_out = 24'b000000000000011100101100;
    16'b1111101000000110 : data_out = 24'b000000000000011100101110;
    16'b1111101000000111 : data_out = 24'b000000000000011100110000;
    16'b1111101000001000 : data_out = 24'b000000000000011100110010;
    16'b1111101000001001 : data_out = 24'b000000000000011100110100;
    16'b1111101000001010 : data_out = 24'b000000000000011100110101;
    16'b1111101000001011 : data_out = 24'b000000000000011100110111;
    16'b1111101000001100 : data_out = 24'b000000000000011100111001;
    16'b1111101000001101 : data_out = 24'b000000000000011100111011;
    16'b1111101000001110 : data_out = 24'b000000000000011100111101;
    16'b1111101000001111 : data_out = 24'b000000000000011100111110;
    16'b1111101000010000 : data_out = 24'b000000000000011101000000;
    16'b1111101000010001 : data_out = 24'b000000000000011101000010;
    16'b1111101000010010 : data_out = 24'b000000000000011101000100;
    16'b1111101000010011 : data_out = 24'b000000000000011101000110;
    16'b1111101000010100 : data_out = 24'b000000000000011101000111;
    16'b1111101000010101 : data_out = 24'b000000000000011101001001;
    16'b1111101000010110 : data_out = 24'b000000000000011101001011;
    16'b1111101000010111 : data_out = 24'b000000000000011101001101;
    16'b1111101000011000 : data_out = 24'b000000000000011101001111;
    16'b1111101000011001 : data_out = 24'b000000000000011101010001;
    16'b1111101000011010 : data_out = 24'b000000000000011101010010;
    16'b1111101000011011 : data_out = 24'b000000000000011101010100;
    16'b1111101000011100 : data_out = 24'b000000000000011101010110;
    16'b1111101000011101 : data_out = 24'b000000000000011101011000;
    16'b1111101000011110 : data_out = 24'b000000000000011101011010;
    16'b1111101000011111 : data_out = 24'b000000000000011101011100;
    16'b1111101000100000 : data_out = 24'b000000000000011101011101;
    16'b1111101000100001 : data_out = 24'b000000000000011101011111;
    16'b1111101000100010 : data_out = 24'b000000000000011101100001;
    16'b1111101000100011 : data_out = 24'b000000000000011101100011;
    16'b1111101000100100 : data_out = 24'b000000000000011101100101;
    16'b1111101000100101 : data_out = 24'b000000000000011101100111;
    16'b1111101000100110 : data_out = 24'b000000000000011101101000;
    16'b1111101000100111 : data_out = 24'b000000000000011101101010;
    16'b1111101000101000 : data_out = 24'b000000000000011101101100;
    16'b1111101000101001 : data_out = 24'b000000000000011101101110;
    16'b1111101000101010 : data_out = 24'b000000000000011101110000;
    16'b1111101000101011 : data_out = 24'b000000000000011101110010;
    16'b1111101000101100 : data_out = 24'b000000000000011101110100;
    16'b1111101000101101 : data_out = 24'b000000000000011101110110;
    16'b1111101000101110 : data_out = 24'b000000000000011101110111;
    16'b1111101000101111 : data_out = 24'b000000000000011101111001;
    16'b1111101000110000 : data_out = 24'b000000000000011101111011;
    16'b1111101000110001 : data_out = 24'b000000000000011101111101;
    16'b1111101000110010 : data_out = 24'b000000000000011101111111;
    16'b1111101000110011 : data_out = 24'b000000000000011110000001;
    16'b1111101000110100 : data_out = 24'b000000000000011110000011;
    16'b1111101000110101 : data_out = 24'b000000000000011110000100;
    16'b1111101000110110 : data_out = 24'b000000000000011110000110;
    16'b1111101000110111 : data_out = 24'b000000000000011110001000;
    16'b1111101000111000 : data_out = 24'b000000000000011110001010;
    16'b1111101000111001 : data_out = 24'b000000000000011110001100;
    16'b1111101000111010 : data_out = 24'b000000000000011110001110;
    16'b1111101000111011 : data_out = 24'b000000000000011110010000;
    16'b1111101000111100 : data_out = 24'b000000000000011110010010;
    16'b1111101000111101 : data_out = 24'b000000000000011110010100;
    16'b1111101000111110 : data_out = 24'b000000000000011110010101;
    16'b1111101000111111 : data_out = 24'b000000000000011110010111;
    16'b1111101001000000 : data_out = 24'b000000000000011110011001;
    16'b1111101001000001 : data_out = 24'b000000000000011110011011;
    16'b1111101001000010 : data_out = 24'b000000000000011110011101;
    16'b1111101001000011 : data_out = 24'b000000000000011110011111;
    16'b1111101001000100 : data_out = 24'b000000000000011110100001;
    16'b1111101001000101 : data_out = 24'b000000000000011110100011;
    16'b1111101001000110 : data_out = 24'b000000000000011110100101;
    16'b1111101001000111 : data_out = 24'b000000000000011110100111;
    16'b1111101001001000 : data_out = 24'b000000000000011110101001;
    16'b1111101001001001 : data_out = 24'b000000000000011110101010;
    16'b1111101001001010 : data_out = 24'b000000000000011110101100;
    16'b1111101001001011 : data_out = 24'b000000000000011110101110;
    16'b1111101001001100 : data_out = 24'b000000000000011110110000;
    16'b1111101001001101 : data_out = 24'b000000000000011110110010;
    16'b1111101001001110 : data_out = 24'b000000000000011110110100;
    16'b1111101001001111 : data_out = 24'b000000000000011110110110;
    16'b1111101001010000 : data_out = 24'b000000000000011110111000;
    16'b1111101001010001 : data_out = 24'b000000000000011110111010;
    16'b1111101001010010 : data_out = 24'b000000000000011110111100;
    16'b1111101001010011 : data_out = 24'b000000000000011110111110;
    16'b1111101001010100 : data_out = 24'b000000000000011111000000;
    16'b1111101001010101 : data_out = 24'b000000000000011111000010;
    16'b1111101001010110 : data_out = 24'b000000000000011111000100;
    16'b1111101001010111 : data_out = 24'b000000000000011111000101;
    16'b1111101001011000 : data_out = 24'b000000000000011111000111;
    16'b1111101001011001 : data_out = 24'b000000000000011111001001;
    16'b1111101001011010 : data_out = 24'b000000000000011111001011;
    16'b1111101001011011 : data_out = 24'b000000000000011111001101;
    16'b1111101001011100 : data_out = 24'b000000000000011111001111;
    16'b1111101001011101 : data_out = 24'b000000000000011111010001;
    16'b1111101001011110 : data_out = 24'b000000000000011111010011;
    16'b1111101001011111 : data_out = 24'b000000000000011111010101;
    16'b1111101001100000 : data_out = 24'b000000000000011111010111;
    16'b1111101001100001 : data_out = 24'b000000000000011111011001;
    16'b1111101001100010 : data_out = 24'b000000000000011111011011;
    16'b1111101001100011 : data_out = 24'b000000000000011111011101;
    16'b1111101001100100 : data_out = 24'b000000000000011111011111;
    16'b1111101001100101 : data_out = 24'b000000000000011111100001;
    16'b1111101001100110 : data_out = 24'b000000000000011111100011;
    16'b1111101001100111 : data_out = 24'b000000000000011111100101;
    16'b1111101001101000 : data_out = 24'b000000000000011111100111;
    16'b1111101001101001 : data_out = 24'b000000000000011111101001;
    16'b1111101001101010 : data_out = 24'b000000000000011111101011;
    16'b1111101001101011 : data_out = 24'b000000000000011111101101;
    16'b1111101001101100 : data_out = 24'b000000000000011111101111;
    16'b1111101001101101 : data_out = 24'b000000000000011111110001;
    16'b1111101001101110 : data_out = 24'b000000000000011111110011;
    16'b1111101001101111 : data_out = 24'b000000000000011111110101;
    16'b1111101001110000 : data_out = 24'b000000000000011111110111;
    16'b1111101001110001 : data_out = 24'b000000000000011111111001;
    16'b1111101001110010 : data_out = 24'b000000000000011111111011;
    16'b1111101001110011 : data_out = 24'b000000000000011111111101;
    16'b1111101001110100 : data_out = 24'b000000000000011111111111;
    16'b1111101001110101 : data_out = 24'b000000000000100000000001;
    16'b1111101001110110 : data_out = 24'b000000000000100000000011;
    16'b1111101001110111 : data_out = 24'b000000000000100000000101;
    16'b1111101001111000 : data_out = 24'b000000000000100000000111;
    16'b1111101001111001 : data_out = 24'b000000000000100000001001;
    16'b1111101001111010 : data_out = 24'b000000000000100000001011;
    16'b1111101001111011 : data_out = 24'b000000000000100000001101;
    16'b1111101001111100 : data_out = 24'b000000000000100000001111;
    16'b1111101001111101 : data_out = 24'b000000000000100000010001;
    16'b1111101001111110 : data_out = 24'b000000000000100000010011;
    16'b1111101001111111 : data_out = 24'b000000000000100000010101;
    16'b1111101010000000 : data_out = 24'b000000000000100000010111;
    16'b1111101010000001 : data_out = 24'b000000000000100000011001;
    16'b1111101010000010 : data_out = 24'b000000000000100000011011;
    16'b1111101010000011 : data_out = 24'b000000000000100000011101;
    16'b1111101010000100 : data_out = 24'b000000000000100000011111;
    16'b1111101010000101 : data_out = 24'b000000000000100000100001;
    16'b1111101010000110 : data_out = 24'b000000000000100000100011;
    16'b1111101010000111 : data_out = 24'b000000000000100000100101;
    16'b1111101010001000 : data_out = 24'b000000000000100000100111;
    16'b1111101010001001 : data_out = 24'b000000000000100000101001;
    16'b1111101010001010 : data_out = 24'b000000000000100000101011;
    16'b1111101010001011 : data_out = 24'b000000000000100000101101;
    16'b1111101010001100 : data_out = 24'b000000000000100000101111;
    16'b1111101010001101 : data_out = 24'b000000000000100000110001;
    16'b1111101010001110 : data_out = 24'b000000000000100000110011;
    16'b1111101010001111 : data_out = 24'b000000000000100000110101;
    16'b1111101010010000 : data_out = 24'b000000000000100000110111;
    16'b1111101010010001 : data_out = 24'b000000000000100000111001;
    16'b1111101010010010 : data_out = 24'b000000000000100000111011;
    16'b1111101010010011 : data_out = 24'b000000000000100000111110;
    16'b1111101010010100 : data_out = 24'b000000000000100001000000;
    16'b1111101010010101 : data_out = 24'b000000000000100001000010;
    16'b1111101010010110 : data_out = 24'b000000000000100001000100;
    16'b1111101010010111 : data_out = 24'b000000000000100001000110;
    16'b1111101010011000 : data_out = 24'b000000000000100001001000;
    16'b1111101010011001 : data_out = 24'b000000000000100001001010;
    16'b1111101010011010 : data_out = 24'b000000000000100001001100;
    16'b1111101010011011 : data_out = 24'b000000000000100001001110;
    16'b1111101010011100 : data_out = 24'b000000000000100001010000;
    16'b1111101010011101 : data_out = 24'b000000000000100001010010;
    16'b1111101010011110 : data_out = 24'b000000000000100001010100;
    16'b1111101010011111 : data_out = 24'b000000000000100001010110;
    16'b1111101010100000 : data_out = 24'b000000000000100001011001;
    16'b1111101010100001 : data_out = 24'b000000000000100001011011;
    16'b1111101010100010 : data_out = 24'b000000000000100001011101;
    16'b1111101010100011 : data_out = 24'b000000000000100001011111;
    16'b1111101010100100 : data_out = 24'b000000000000100001100001;
    16'b1111101010100101 : data_out = 24'b000000000000100001100011;
    16'b1111101010100110 : data_out = 24'b000000000000100001100101;
    16'b1111101010100111 : data_out = 24'b000000000000100001100111;
    16'b1111101010101000 : data_out = 24'b000000000000100001101001;
    16'b1111101010101001 : data_out = 24'b000000000000100001101011;
    16'b1111101010101010 : data_out = 24'b000000000000100001101101;
    16'b1111101010101011 : data_out = 24'b000000000000100001110000;
    16'b1111101010101100 : data_out = 24'b000000000000100001110010;
    16'b1111101010101101 : data_out = 24'b000000000000100001110100;
    16'b1111101010101110 : data_out = 24'b000000000000100001110110;
    16'b1111101010101111 : data_out = 24'b000000000000100001111000;
    16'b1111101010110000 : data_out = 24'b000000000000100001111010;
    16'b1111101010110001 : data_out = 24'b000000000000100001111100;
    16'b1111101010110010 : data_out = 24'b000000000000100001111110;
    16'b1111101010110011 : data_out = 24'b000000000000100010000001;
    16'b1111101010110100 : data_out = 24'b000000000000100010000011;
    16'b1111101010110101 : data_out = 24'b000000000000100010000101;
    16'b1111101010110110 : data_out = 24'b000000000000100010000111;
    16'b1111101010110111 : data_out = 24'b000000000000100010001001;
    16'b1111101010111000 : data_out = 24'b000000000000100010001011;
    16'b1111101010111001 : data_out = 24'b000000000000100010001101;
    16'b1111101010111010 : data_out = 24'b000000000000100010001111;
    16'b1111101010111011 : data_out = 24'b000000000000100010010010;
    16'b1111101010111100 : data_out = 24'b000000000000100010010100;
    16'b1111101010111101 : data_out = 24'b000000000000100010010110;
    16'b1111101010111110 : data_out = 24'b000000000000100010011000;
    16'b1111101010111111 : data_out = 24'b000000000000100010011010;
    16'b1111101011000000 : data_out = 24'b000000000000100010011100;
    16'b1111101011000001 : data_out = 24'b000000000000100010011111;
    16'b1111101011000010 : data_out = 24'b000000000000100010100001;
    16'b1111101011000011 : data_out = 24'b000000000000100010100011;
    16'b1111101011000100 : data_out = 24'b000000000000100010100101;
    16'b1111101011000101 : data_out = 24'b000000000000100010100111;
    16'b1111101011000110 : data_out = 24'b000000000000100010101001;
    16'b1111101011000111 : data_out = 24'b000000000000100010101011;
    16'b1111101011001000 : data_out = 24'b000000000000100010101110;
    16'b1111101011001001 : data_out = 24'b000000000000100010110000;
    16'b1111101011001010 : data_out = 24'b000000000000100010110010;
    16'b1111101011001011 : data_out = 24'b000000000000100010110100;
    16'b1111101011001100 : data_out = 24'b000000000000100010110110;
    16'b1111101011001101 : data_out = 24'b000000000000100010111001;
    16'b1111101011001110 : data_out = 24'b000000000000100010111011;
    16'b1111101011001111 : data_out = 24'b000000000000100010111101;
    16'b1111101011010000 : data_out = 24'b000000000000100010111111;
    16'b1111101011010001 : data_out = 24'b000000000000100011000001;
    16'b1111101011010010 : data_out = 24'b000000000000100011000011;
    16'b1111101011010011 : data_out = 24'b000000000000100011000110;
    16'b1111101011010100 : data_out = 24'b000000000000100011001000;
    16'b1111101011010101 : data_out = 24'b000000000000100011001010;
    16'b1111101011010110 : data_out = 24'b000000000000100011001100;
    16'b1111101011010111 : data_out = 24'b000000000000100011001110;
    16'b1111101011011000 : data_out = 24'b000000000000100011010001;
    16'b1111101011011001 : data_out = 24'b000000000000100011010011;
    16'b1111101011011010 : data_out = 24'b000000000000100011010101;
    16'b1111101011011011 : data_out = 24'b000000000000100011010111;
    16'b1111101011011100 : data_out = 24'b000000000000100011011001;
    16'b1111101011011101 : data_out = 24'b000000000000100011011100;
    16'b1111101011011110 : data_out = 24'b000000000000100011011110;
    16'b1111101011011111 : data_out = 24'b000000000000100011100000;
    16'b1111101011100000 : data_out = 24'b000000000000100011100010;
    16'b1111101011100001 : data_out = 24'b000000000000100011100101;
    16'b1111101011100010 : data_out = 24'b000000000000100011100111;
    16'b1111101011100011 : data_out = 24'b000000000000100011101001;
    16'b1111101011100100 : data_out = 24'b000000000000100011101011;
    16'b1111101011100101 : data_out = 24'b000000000000100011101101;
    16'b1111101011100110 : data_out = 24'b000000000000100011110000;
    16'b1111101011100111 : data_out = 24'b000000000000100011110010;
    16'b1111101011101000 : data_out = 24'b000000000000100011110100;
    16'b1111101011101001 : data_out = 24'b000000000000100011110110;
    16'b1111101011101010 : data_out = 24'b000000000000100011111001;
    16'b1111101011101011 : data_out = 24'b000000000000100011111011;
    16'b1111101011101100 : data_out = 24'b000000000000100011111101;
    16'b1111101011101101 : data_out = 24'b000000000000100011111111;
    16'b1111101011101110 : data_out = 24'b000000000000100100000010;
    16'b1111101011101111 : data_out = 24'b000000000000100100000100;
    16'b1111101011110000 : data_out = 24'b000000000000100100000110;
    16'b1111101011110001 : data_out = 24'b000000000000100100001000;
    16'b1111101011110010 : data_out = 24'b000000000000100100001011;
    16'b1111101011110011 : data_out = 24'b000000000000100100001101;
    16'b1111101011110100 : data_out = 24'b000000000000100100001111;
    16'b1111101011110101 : data_out = 24'b000000000000100100010001;
    16'b1111101011110110 : data_out = 24'b000000000000100100010100;
    16'b1111101011110111 : data_out = 24'b000000000000100100010110;
    16'b1111101011111000 : data_out = 24'b000000000000100100011000;
    16'b1111101011111001 : data_out = 24'b000000000000100100011011;
    16'b1111101011111010 : data_out = 24'b000000000000100100011101;
    16'b1111101011111011 : data_out = 24'b000000000000100100011111;
    16'b1111101011111100 : data_out = 24'b000000000000100100100001;
    16'b1111101011111101 : data_out = 24'b000000000000100100100100;
    16'b1111101011111110 : data_out = 24'b000000000000100100100110;
    16'b1111101011111111 : data_out = 24'b000000000000100100101000;
    16'b1111101100000000 : data_out = 24'b000000000000100100101011;
    16'b1111101100000001 : data_out = 24'b000000000000100100101101;
    16'b1111101100000010 : data_out = 24'b000000000000100100101111;
    16'b1111101100000011 : data_out = 24'b000000000000100100110001;
    16'b1111101100000100 : data_out = 24'b000000000000100100110100;
    16'b1111101100000101 : data_out = 24'b000000000000100100110110;
    16'b1111101100000110 : data_out = 24'b000000000000100100111000;
    16'b1111101100000111 : data_out = 24'b000000000000100100111011;
    16'b1111101100001000 : data_out = 24'b000000000000100100111101;
    16'b1111101100001001 : data_out = 24'b000000000000100100111111;
    16'b1111101100001010 : data_out = 24'b000000000000100101000010;
    16'b1111101100001011 : data_out = 24'b000000000000100101000100;
    16'b1111101100001100 : data_out = 24'b000000000000100101000110;
    16'b1111101100001101 : data_out = 24'b000000000000100101001001;
    16'b1111101100001110 : data_out = 24'b000000000000100101001011;
    16'b1111101100001111 : data_out = 24'b000000000000100101001101;
    16'b1111101100010000 : data_out = 24'b000000000000100101010000;
    16'b1111101100010001 : data_out = 24'b000000000000100101010010;
    16'b1111101100010010 : data_out = 24'b000000000000100101010100;
    16'b1111101100010011 : data_out = 24'b000000000000100101010111;
    16'b1111101100010100 : data_out = 24'b000000000000100101011001;
    16'b1111101100010101 : data_out = 24'b000000000000100101011011;
    16'b1111101100010110 : data_out = 24'b000000000000100101011110;
    16'b1111101100010111 : data_out = 24'b000000000000100101100000;
    16'b1111101100011000 : data_out = 24'b000000000000100101100010;
    16'b1111101100011001 : data_out = 24'b000000000000100101100101;
    16'b1111101100011010 : data_out = 24'b000000000000100101100111;
    16'b1111101100011011 : data_out = 24'b000000000000100101101001;
    16'b1111101100011100 : data_out = 24'b000000000000100101101100;
    16'b1111101100011101 : data_out = 24'b000000000000100101101110;
    16'b1111101100011110 : data_out = 24'b000000000000100101110000;
    16'b1111101100011111 : data_out = 24'b000000000000100101110011;
    16'b1111101100100000 : data_out = 24'b000000000000100101110101;
    16'b1111101100100001 : data_out = 24'b000000000000100101110111;
    16'b1111101100100010 : data_out = 24'b000000000000100101111010;
    16'b1111101100100011 : data_out = 24'b000000000000100101111100;
    16'b1111101100100100 : data_out = 24'b000000000000100101111111;
    16'b1111101100100101 : data_out = 24'b000000000000100110000001;
    16'b1111101100100110 : data_out = 24'b000000000000100110000011;
    16'b1111101100100111 : data_out = 24'b000000000000100110000110;
    16'b1111101100101000 : data_out = 24'b000000000000100110001000;
    16'b1111101100101001 : data_out = 24'b000000000000100110001010;
    16'b1111101100101010 : data_out = 24'b000000000000100110001101;
    16'b1111101100101011 : data_out = 24'b000000000000100110001111;
    16'b1111101100101100 : data_out = 24'b000000000000100110010010;
    16'b1111101100101101 : data_out = 24'b000000000000100110010100;
    16'b1111101100101110 : data_out = 24'b000000000000100110010110;
    16'b1111101100101111 : data_out = 24'b000000000000100110011001;
    16'b1111101100110000 : data_out = 24'b000000000000100110011011;
    16'b1111101100110001 : data_out = 24'b000000000000100110011110;
    16'b1111101100110010 : data_out = 24'b000000000000100110100000;
    16'b1111101100110011 : data_out = 24'b000000000000100110100010;
    16'b1111101100110100 : data_out = 24'b000000000000100110100101;
    16'b1111101100110101 : data_out = 24'b000000000000100110100111;
    16'b1111101100110110 : data_out = 24'b000000000000100110101010;
    16'b1111101100110111 : data_out = 24'b000000000000100110101100;
    16'b1111101100111000 : data_out = 24'b000000000000100110101110;
    16'b1111101100111001 : data_out = 24'b000000000000100110110001;
    16'b1111101100111010 : data_out = 24'b000000000000100110110011;
    16'b1111101100111011 : data_out = 24'b000000000000100110110110;
    16'b1111101100111100 : data_out = 24'b000000000000100110111000;
    16'b1111101100111101 : data_out = 24'b000000000000100110111011;
    16'b1111101100111110 : data_out = 24'b000000000000100110111101;
    16'b1111101100111111 : data_out = 24'b000000000000100110111111;
    16'b1111101101000000 : data_out = 24'b000000000000100111000010;
    16'b1111101101000001 : data_out = 24'b000000000000100111000100;
    16'b1111101101000010 : data_out = 24'b000000000000100111000111;
    16'b1111101101000011 : data_out = 24'b000000000000100111001001;
    16'b1111101101000100 : data_out = 24'b000000000000100111001100;
    16'b1111101101000101 : data_out = 24'b000000000000100111001110;
    16'b1111101101000110 : data_out = 24'b000000000000100111010001;
    16'b1111101101000111 : data_out = 24'b000000000000100111010011;
    16'b1111101101001000 : data_out = 24'b000000000000100111010110;
    16'b1111101101001001 : data_out = 24'b000000000000100111011000;
    16'b1111101101001010 : data_out = 24'b000000000000100111011010;
    16'b1111101101001011 : data_out = 24'b000000000000100111011101;
    16'b1111101101001100 : data_out = 24'b000000000000100111011111;
    16'b1111101101001101 : data_out = 24'b000000000000100111100010;
    16'b1111101101001110 : data_out = 24'b000000000000100111100100;
    16'b1111101101001111 : data_out = 24'b000000000000100111100111;
    16'b1111101101010000 : data_out = 24'b000000000000100111101001;
    16'b1111101101010001 : data_out = 24'b000000000000100111101100;
    16'b1111101101010010 : data_out = 24'b000000000000100111101110;
    16'b1111101101010011 : data_out = 24'b000000000000100111110001;
    16'b1111101101010100 : data_out = 24'b000000000000100111110011;
    16'b1111101101010101 : data_out = 24'b000000000000100111110110;
    16'b1111101101010110 : data_out = 24'b000000000000100111111000;
    16'b1111101101010111 : data_out = 24'b000000000000100111111011;
    16'b1111101101011000 : data_out = 24'b000000000000100111111101;
    16'b1111101101011001 : data_out = 24'b000000000000101000000000;
    16'b1111101101011010 : data_out = 24'b000000000000101000000010;
    16'b1111101101011011 : data_out = 24'b000000000000101000000101;
    16'b1111101101011100 : data_out = 24'b000000000000101000000111;
    16'b1111101101011101 : data_out = 24'b000000000000101000001010;
    16'b1111101101011110 : data_out = 24'b000000000000101000001100;
    16'b1111101101011111 : data_out = 24'b000000000000101000001111;
    16'b1111101101100000 : data_out = 24'b000000000000101000010001;
    16'b1111101101100001 : data_out = 24'b000000000000101000010100;
    16'b1111101101100010 : data_out = 24'b000000000000101000010110;
    16'b1111101101100011 : data_out = 24'b000000000000101000011001;
    16'b1111101101100100 : data_out = 24'b000000000000101000011011;
    16'b1111101101100101 : data_out = 24'b000000000000101000011110;
    16'b1111101101100110 : data_out = 24'b000000000000101000100000;
    16'b1111101101100111 : data_out = 24'b000000000000101000100011;
    16'b1111101101101000 : data_out = 24'b000000000000101000100101;
    16'b1111101101101001 : data_out = 24'b000000000000101000101000;
    16'b1111101101101010 : data_out = 24'b000000000000101000101011;
    16'b1111101101101011 : data_out = 24'b000000000000101000101101;
    16'b1111101101101100 : data_out = 24'b000000000000101000110000;
    16'b1111101101101101 : data_out = 24'b000000000000101000110010;
    16'b1111101101101110 : data_out = 24'b000000000000101000110101;
    16'b1111101101101111 : data_out = 24'b000000000000101000110111;
    16'b1111101101110000 : data_out = 24'b000000000000101000111010;
    16'b1111101101110001 : data_out = 24'b000000000000101000111100;
    16'b1111101101110010 : data_out = 24'b000000000000101000111111;
    16'b1111101101110011 : data_out = 24'b000000000000101001000010;
    16'b1111101101110100 : data_out = 24'b000000000000101001000100;
    16'b1111101101110101 : data_out = 24'b000000000000101001000111;
    16'b1111101101110110 : data_out = 24'b000000000000101001001001;
    16'b1111101101110111 : data_out = 24'b000000000000101001001100;
    16'b1111101101111000 : data_out = 24'b000000000000101001001110;
    16'b1111101101111001 : data_out = 24'b000000000000101001010001;
    16'b1111101101111010 : data_out = 24'b000000000000101001010100;
    16'b1111101101111011 : data_out = 24'b000000000000101001010110;
    16'b1111101101111100 : data_out = 24'b000000000000101001011001;
    16'b1111101101111101 : data_out = 24'b000000000000101001011011;
    16'b1111101101111110 : data_out = 24'b000000000000101001011110;
    16'b1111101101111111 : data_out = 24'b000000000000101001100000;
    16'b1111101110000000 : data_out = 24'b000000000000101001100011;
    16'b1111101110000001 : data_out = 24'b000000000000101001100110;
    16'b1111101110000010 : data_out = 24'b000000000000101001101000;
    16'b1111101110000011 : data_out = 24'b000000000000101001101011;
    16'b1111101110000100 : data_out = 24'b000000000000101001101101;
    16'b1111101110000101 : data_out = 24'b000000000000101001110000;
    16'b1111101110000110 : data_out = 24'b000000000000101001110011;
    16'b1111101110000111 : data_out = 24'b000000000000101001110101;
    16'b1111101110001000 : data_out = 24'b000000000000101001111000;
    16'b1111101110001001 : data_out = 24'b000000000000101001111011;
    16'b1111101110001010 : data_out = 24'b000000000000101001111101;
    16'b1111101110001011 : data_out = 24'b000000000000101010000000;
    16'b1111101110001100 : data_out = 24'b000000000000101010000010;
    16'b1111101110001101 : data_out = 24'b000000000000101010000101;
    16'b1111101110001110 : data_out = 24'b000000000000101010001000;
    16'b1111101110001111 : data_out = 24'b000000000000101010001010;
    16'b1111101110010000 : data_out = 24'b000000000000101010001101;
    16'b1111101110010001 : data_out = 24'b000000000000101010010000;
    16'b1111101110010010 : data_out = 24'b000000000000101010010010;
    16'b1111101110010011 : data_out = 24'b000000000000101010010101;
    16'b1111101110010100 : data_out = 24'b000000000000101010011000;
    16'b1111101110010101 : data_out = 24'b000000000000101010011010;
    16'b1111101110010110 : data_out = 24'b000000000000101010011101;
    16'b1111101110010111 : data_out = 24'b000000000000101010011111;
    16'b1111101110011000 : data_out = 24'b000000000000101010100010;
    16'b1111101110011001 : data_out = 24'b000000000000101010100101;
    16'b1111101110011010 : data_out = 24'b000000000000101010100111;
    16'b1111101110011011 : data_out = 24'b000000000000101010101010;
    16'b1111101110011100 : data_out = 24'b000000000000101010101101;
    16'b1111101110011101 : data_out = 24'b000000000000101010101111;
    16'b1111101110011110 : data_out = 24'b000000000000101010110010;
    16'b1111101110011111 : data_out = 24'b000000000000101010110101;
    16'b1111101110100000 : data_out = 24'b000000000000101010110111;
    16'b1111101110100001 : data_out = 24'b000000000000101010111010;
    16'b1111101110100010 : data_out = 24'b000000000000101010111101;
    16'b1111101110100011 : data_out = 24'b000000000000101011000000;
    16'b1111101110100100 : data_out = 24'b000000000000101011000010;
    16'b1111101110100101 : data_out = 24'b000000000000101011000101;
    16'b1111101110100110 : data_out = 24'b000000000000101011001000;
    16'b1111101110100111 : data_out = 24'b000000000000101011001010;
    16'b1111101110101000 : data_out = 24'b000000000000101011001101;
    16'b1111101110101001 : data_out = 24'b000000000000101011010000;
    16'b1111101110101010 : data_out = 24'b000000000000101011010010;
    16'b1111101110101011 : data_out = 24'b000000000000101011010101;
    16'b1111101110101100 : data_out = 24'b000000000000101011011000;
    16'b1111101110101101 : data_out = 24'b000000000000101011011011;
    16'b1111101110101110 : data_out = 24'b000000000000101011011101;
    16'b1111101110101111 : data_out = 24'b000000000000101011100000;
    16'b1111101110110000 : data_out = 24'b000000000000101011100011;
    16'b1111101110110001 : data_out = 24'b000000000000101011100101;
    16'b1111101110110010 : data_out = 24'b000000000000101011101000;
    16'b1111101110110011 : data_out = 24'b000000000000101011101011;
    16'b1111101110110100 : data_out = 24'b000000000000101011101110;
    16'b1111101110110101 : data_out = 24'b000000000000101011110000;
    16'b1111101110110110 : data_out = 24'b000000000000101011110011;
    16'b1111101110110111 : data_out = 24'b000000000000101011110110;
    16'b1111101110111000 : data_out = 24'b000000000000101011111001;
    16'b1111101110111001 : data_out = 24'b000000000000101011111011;
    16'b1111101110111010 : data_out = 24'b000000000000101011111110;
    16'b1111101110111011 : data_out = 24'b000000000000101100000001;
    16'b1111101110111100 : data_out = 24'b000000000000101100000100;
    16'b1111101110111101 : data_out = 24'b000000000000101100000110;
    16'b1111101110111110 : data_out = 24'b000000000000101100001001;
    16'b1111101110111111 : data_out = 24'b000000000000101100001100;
    16'b1111101111000000 : data_out = 24'b000000000000101100001111;
    16'b1111101111000001 : data_out = 24'b000000000000101100010001;
    16'b1111101111000010 : data_out = 24'b000000000000101100010100;
    16'b1111101111000011 : data_out = 24'b000000000000101100010111;
    16'b1111101111000100 : data_out = 24'b000000000000101100011010;
    16'b1111101111000101 : data_out = 24'b000000000000101100011100;
    16'b1111101111000110 : data_out = 24'b000000000000101100011111;
    16'b1111101111000111 : data_out = 24'b000000000000101100100010;
    16'b1111101111001000 : data_out = 24'b000000000000101100100101;
    16'b1111101111001001 : data_out = 24'b000000000000101100101000;
    16'b1111101111001010 : data_out = 24'b000000000000101100101010;
    16'b1111101111001011 : data_out = 24'b000000000000101100101101;
    16'b1111101111001100 : data_out = 24'b000000000000101100110000;
    16'b1111101111001101 : data_out = 24'b000000000000101100110011;
    16'b1111101111001110 : data_out = 24'b000000000000101100110110;
    16'b1111101111001111 : data_out = 24'b000000000000101100111000;
    16'b1111101111010000 : data_out = 24'b000000000000101100111011;
    16'b1111101111010001 : data_out = 24'b000000000000101100111110;
    16'b1111101111010010 : data_out = 24'b000000000000101101000001;
    16'b1111101111010011 : data_out = 24'b000000000000101101000100;
    16'b1111101111010100 : data_out = 24'b000000000000101101000110;
    16'b1111101111010101 : data_out = 24'b000000000000101101001001;
    16'b1111101111010110 : data_out = 24'b000000000000101101001100;
    16'b1111101111010111 : data_out = 24'b000000000000101101001111;
    16'b1111101111011000 : data_out = 24'b000000000000101101010010;
    16'b1111101111011001 : data_out = 24'b000000000000101101010101;
    16'b1111101111011010 : data_out = 24'b000000000000101101010111;
    16'b1111101111011011 : data_out = 24'b000000000000101101011010;
    16'b1111101111011100 : data_out = 24'b000000000000101101011101;
    16'b1111101111011101 : data_out = 24'b000000000000101101100000;
    16'b1111101111011110 : data_out = 24'b000000000000101101100011;
    16'b1111101111011111 : data_out = 24'b000000000000101101100110;
    16'b1111101111100000 : data_out = 24'b000000000000101101101000;
    16'b1111101111100001 : data_out = 24'b000000000000101101101011;
    16'b1111101111100010 : data_out = 24'b000000000000101101101110;
    16'b1111101111100011 : data_out = 24'b000000000000101101110001;
    16'b1111101111100100 : data_out = 24'b000000000000101101110100;
    16'b1111101111100101 : data_out = 24'b000000000000101101110111;
    16'b1111101111100110 : data_out = 24'b000000000000101101111010;
    16'b1111101111100111 : data_out = 24'b000000000000101101111100;
    16'b1111101111101000 : data_out = 24'b000000000000101101111111;
    16'b1111101111101001 : data_out = 24'b000000000000101110000010;
    16'b1111101111101010 : data_out = 24'b000000000000101110000101;
    16'b1111101111101011 : data_out = 24'b000000000000101110001000;
    16'b1111101111101100 : data_out = 24'b000000000000101110001011;
    16'b1111101111101101 : data_out = 24'b000000000000101110001110;
    16'b1111101111101110 : data_out = 24'b000000000000101110010001;
    16'b1111101111101111 : data_out = 24'b000000000000101110010100;
    16'b1111101111110000 : data_out = 24'b000000000000101110010110;
    16'b1111101111110001 : data_out = 24'b000000000000101110011001;
    16'b1111101111110010 : data_out = 24'b000000000000101110011100;
    16'b1111101111110011 : data_out = 24'b000000000000101110011111;
    16'b1111101111110100 : data_out = 24'b000000000000101110100010;
    16'b1111101111110101 : data_out = 24'b000000000000101110100101;
    16'b1111101111110110 : data_out = 24'b000000000000101110101000;
    16'b1111101111110111 : data_out = 24'b000000000000101110101011;
    16'b1111101111111000 : data_out = 24'b000000000000101110101110;
    16'b1111101111111001 : data_out = 24'b000000000000101110110001;
    16'b1111101111111010 : data_out = 24'b000000000000101110110100;
    16'b1111101111111011 : data_out = 24'b000000000000101110110110;
    16'b1111101111111100 : data_out = 24'b000000000000101110111001;
    16'b1111101111111101 : data_out = 24'b000000000000101110111100;
    16'b1111101111111110 : data_out = 24'b000000000000101110111111;
    16'b1111101111111111 : data_out = 24'b000000000000101111000010;
    16'b1111110000000000 : data_out = 24'b000000000000101111000101;
    16'b1111110000000001 : data_out = 24'b000000000000101111001000;
    16'b1111110000000010 : data_out = 24'b000000000000101111001011;
    16'b1111110000000011 : data_out = 24'b000000000000101111001110;
    16'b1111110000000100 : data_out = 24'b000000000000101111010001;
    16'b1111110000000101 : data_out = 24'b000000000000101111010100;
    16'b1111110000000110 : data_out = 24'b000000000000101111010111;
    16'b1111110000000111 : data_out = 24'b000000000000101111011010;
    16'b1111110000001000 : data_out = 24'b000000000000101111011101;
    16'b1111110000001001 : data_out = 24'b000000000000101111100000;
    16'b1111110000001010 : data_out = 24'b000000000000101111100011;
    16'b1111110000001011 : data_out = 24'b000000000000101111100110;
    16'b1111110000001100 : data_out = 24'b000000000000101111101001;
    16'b1111110000001101 : data_out = 24'b000000000000101111101100;
    16'b1111110000001110 : data_out = 24'b000000000000101111101111;
    16'b1111110000001111 : data_out = 24'b000000000000101111110010;
    16'b1111110000010000 : data_out = 24'b000000000000101111110101;
    16'b1111110000010001 : data_out = 24'b000000000000101111111000;
    16'b1111110000010010 : data_out = 24'b000000000000101111111011;
    16'b1111110000010011 : data_out = 24'b000000000000101111111110;
    16'b1111110000010100 : data_out = 24'b000000000000110000000001;
    16'b1111110000010101 : data_out = 24'b000000000000110000000100;
    16'b1111110000010110 : data_out = 24'b000000000000110000000111;
    16'b1111110000010111 : data_out = 24'b000000000000110000001010;
    16'b1111110000011000 : data_out = 24'b000000000000110000001101;
    16'b1111110000011001 : data_out = 24'b000000000000110000010000;
    16'b1111110000011010 : data_out = 24'b000000000000110000010011;
    16'b1111110000011011 : data_out = 24'b000000000000110000010110;
    16'b1111110000011100 : data_out = 24'b000000000000110000011001;
    16'b1111110000011101 : data_out = 24'b000000000000110000011100;
    16'b1111110000011110 : data_out = 24'b000000000000110000011111;
    16'b1111110000011111 : data_out = 24'b000000000000110000100010;
    16'b1111110000100000 : data_out = 24'b000000000000110000100101;
    16'b1111110000100001 : data_out = 24'b000000000000110000101000;
    16'b1111110000100010 : data_out = 24'b000000000000110000101011;
    16'b1111110000100011 : data_out = 24'b000000000000110000101110;
    16'b1111110000100100 : data_out = 24'b000000000000110000110001;
    16'b1111110000100101 : data_out = 24'b000000000000110000110100;
    16'b1111110000100110 : data_out = 24'b000000000000110000110111;
    16'b1111110000100111 : data_out = 24'b000000000000110000111010;
    16'b1111110000101000 : data_out = 24'b000000000000110000111101;
    16'b1111110000101001 : data_out = 24'b000000000000110001000000;
    16'b1111110000101010 : data_out = 24'b000000000000110001000011;
    16'b1111110000101011 : data_out = 24'b000000000000110001000110;
    16'b1111110000101100 : data_out = 24'b000000000000110001001001;
    16'b1111110000101101 : data_out = 24'b000000000000110001001101;
    16'b1111110000101110 : data_out = 24'b000000000000110001010000;
    16'b1111110000101111 : data_out = 24'b000000000000110001010011;
    16'b1111110000110000 : data_out = 24'b000000000000110001010110;
    16'b1111110000110001 : data_out = 24'b000000000000110001011001;
    16'b1111110000110010 : data_out = 24'b000000000000110001011100;
    16'b1111110000110011 : data_out = 24'b000000000000110001011111;
    16'b1111110000110100 : data_out = 24'b000000000000110001100010;
    16'b1111110000110101 : data_out = 24'b000000000000110001100101;
    16'b1111110000110110 : data_out = 24'b000000000000110001101000;
    16'b1111110000110111 : data_out = 24'b000000000000110001101011;
    16'b1111110000111000 : data_out = 24'b000000000000110001101111;
    16'b1111110000111001 : data_out = 24'b000000000000110001110010;
    16'b1111110000111010 : data_out = 24'b000000000000110001110101;
    16'b1111110000111011 : data_out = 24'b000000000000110001111000;
    16'b1111110000111100 : data_out = 24'b000000000000110001111011;
    16'b1111110000111101 : data_out = 24'b000000000000110001111110;
    16'b1111110000111110 : data_out = 24'b000000000000110010000001;
    16'b1111110000111111 : data_out = 24'b000000000000110010000100;
    16'b1111110001000000 : data_out = 24'b000000000000110010001000;
    16'b1111110001000001 : data_out = 24'b000000000000110010001011;
    16'b1111110001000010 : data_out = 24'b000000000000110010001110;
    16'b1111110001000011 : data_out = 24'b000000000000110010010001;
    16'b1111110001000100 : data_out = 24'b000000000000110010010100;
    16'b1111110001000101 : data_out = 24'b000000000000110010010111;
    16'b1111110001000110 : data_out = 24'b000000000000110010011010;
    16'b1111110001000111 : data_out = 24'b000000000000110010011110;
    16'b1111110001001000 : data_out = 24'b000000000000110010100001;
    16'b1111110001001001 : data_out = 24'b000000000000110010100100;
    16'b1111110001001010 : data_out = 24'b000000000000110010100111;
    16'b1111110001001011 : data_out = 24'b000000000000110010101010;
    16'b1111110001001100 : data_out = 24'b000000000000110010101101;
    16'b1111110001001101 : data_out = 24'b000000000000110010110001;
    16'b1111110001001110 : data_out = 24'b000000000000110010110100;
    16'b1111110001001111 : data_out = 24'b000000000000110010110111;
    16'b1111110001010000 : data_out = 24'b000000000000110010111010;
    16'b1111110001010001 : data_out = 24'b000000000000110010111101;
    16'b1111110001010010 : data_out = 24'b000000000000110011000000;
    16'b1111110001010011 : data_out = 24'b000000000000110011000100;
    16'b1111110001010100 : data_out = 24'b000000000000110011000111;
    16'b1111110001010101 : data_out = 24'b000000000000110011001010;
    16'b1111110001010110 : data_out = 24'b000000000000110011001101;
    16'b1111110001010111 : data_out = 24'b000000000000110011010000;
    16'b1111110001011000 : data_out = 24'b000000000000110011010100;
    16'b1111110001011001 : data_out = 24'b000000000000110011010111;
    16'b1111110001011010 : data_out = 24'b000000000000110011011010;
    16'b1111110001011011 : data_out = 24'b000000000000110011011101;
    16'b1111110001011100 : data_out = 24'b000000000000110011100000;
    16'b1111110001011101 : data_out = 24'b000000000000110011100100;
    16'b1111110001011110 : data_out = 24'b000000000000110011100111;
    16'b1111110001011111 : data_out = 24'b000000000000110011101010;
    16'b1111110001100000 : data_out = 24'b000000000000110011101101;
    16'b1111110001100001 : data_out = 24'b000000000000110011110001;
    16'b1111110001100010 : data_out = 24'b000000000000110011110100;
    16'b1111110001100011 : data_out = 24'b000000000000110011110111;
    16'b1111110001100100 : data_out = 24'b000000000000110011111010;
    16'b1111110001100101 : data_out = 24'b000000000000110011111110;
    16'b1111110001100110 : data_out = 24'b000000000000110100000001;
    16'b1111110001100111 : data_out = 24'b000000000000110100000100;
    16'b1111110001101000 : data_out = 24'b000000000000110100000111;
    16'b1111110001101001 : data_out = 24'b000000000000110100001011;
    16'b1111110001101010 : data_out = 24'b000000000000110100001110;
    16'b1111110001101011 : data_out = 24'b000000000000110100010001;
    16'b1111110001101100 : data_out = 24'b000000000000110100010100;
    16'b1111110001101101 : data_out = 24'b000000000000110100011000;
    16'b1111110001101110 : data_out = 24'b000000000000110100011011;
    16'b1111110001101111 : data_out = 24'b000000000000110100011110;
    16'b1111110001110000 : data_out = 24'b000000000000110100100001;
    16'b1111110001110001 : data_out = 24'b000000000000110100100101;
    16'b1111110001110010 : data_out = 24'b000000000000110100101000;
    16'b1111110001110011 : data_out = 24'b000000000000110100101011;
    16'b1111110001110100 : data_out = 24'b000000000000110100101111;
    16'b1111110001110101 : data_out = 24'b000000000000110100110010;
    16'b1111110001110110 : data_out = 24'b000000000000110100110101;
    16'b1111110001110111 : data_out = 24'b000000000000110100111001;
    16'b1111110001111000 : data_out = 24'b000000000000110100111100;
    16'b1111110001111001 : data_out = 24'b000000000000110100111111;
    16'b1111110001111010 : data_out = 24'b000000000000110101000010;
    16'b1111110001111011 : data_out = 24'b000000000000110101000110;
    16'b1111110001111100 : data_out = 24'b000000000000110101001001;
    16'b1111110001111101 : data_out = 24'b000000000000110101001100;
    16'b1111110001111110 : data_out = 24'b000000000000110101010000;
    16'b1111110001111111 : data_out = 24'b000000000000110101010011;
    16'b1111110010000000 : data_out = 24'b000000000000110101010110;
    16'b1111110010000001 : data_out = 24'b000000000000110101011010;
    16'b1111110010000010 : data_out = 24'b000000000000110101011101;
    16'b1111110010000011 : data_out = 24'b000000000000110101100000;
    16'b1111110010000100 : data_out = 24'b000000000000110101100100;
    16'b1111110010000101 : data_out = 24'b000000000000110101100111;
    16'b1111110010000110 : data_out = 24'b000000000000110101101011;
    16'b1111110010000111 : data_out = 24'b000000000000110101101110;
    16'b1111110010001000 : data_out = 24'b000000000000110101110001;
    16'b1111110010001001 : data_out = 24'b000000000000110101110101;
    16'b1111110010001010 : data_out = 24'b000000000000110101111000;
    16'b1111110010001011 : data_out = 24'b000000000000110101111011;
    16'b1111110010001100 : data_out = 24'b000000000000110101111111;
    16'b1111110010001101 : data_out = 24'b000000000000110110000010;
    16'b1111110010001110 : data_out = 24'b000000000000110110000101;
    16'b1111110010001111 : data_out = 24'b000000000000110110001001;
    16'b1111110010010000 : data_out = 24'b000000000000110110001100;
    16'b1111110010010001 : data_out = 24'b000000000000110110010000;
    16'b1111110010010010 : data_out = 24'b000000000000110110010011;
    16'b1111110010010011 : data_out = 24'b000000000000110110010110;
    16'b1111110010010100 : data_out = 24'b000000000000110110011010;
    16'b1111110010010101 : data_out = 24'b000000000000110110011101;
    16'b1111110010010110 : data_out = 24'b000000000000110110100001;
    16'b1111110010010111 : data_out = 24'b000000000000110110100100;
    16'b1111110010011000 : data_out = 24'b000000000000110110100111;
    16'b1111110010011001 : data_out = 24'b000000000000110110101011;
    16'b1111110010011010 : data_out = 24'b000000000000110110101110;
    16'b1111110010011011 : data_out = 24'b000000000000110110110010;
    16'b1111110010011100 : data_out = 24'b000000000000110110110101;
    16'b1111110010011101 : data_out = 24'b000000000000110110111001;
    16'b1111110010011110 : data_out = 24'b000000000000110110111100;
    16'b1111110010011111 : data_out = 24'b000000000000110110111111;
    16'b1111110010100000 : data_out = 24'b000000000000110111000011;
    16'b1111110010100001 : data_out = 24'b000000000000110111000110;
    16'b1111110010100010 : data_out = 24'b000000000000110111001010;
    16'b1111110010100011 : data_out = 24'b000000000000110111001101;
    16'b1111110010100100 : data_out = 24'b000000000000110111010001;
    16'b1111110010100101 : data_out = 24'b000000000000110111010100;
    16'b1111110010100110 : data_out = 24'b000000000000110111011000;
    16'b1111110010100111 : data_out = 24'b000000000000110111011011;
    16'b1111110010101000 : data_out = 24'b000000000000110111011110;
    16'b1111110010101001 : data_out = 24'b000000000000110111100010;
    16'b1111110010101010 : data_out = 24'b000000000000110111100101;
    16'b1111110010101011 : data_out = 24'b000000000000110111101001;
    16'b1111110010101100 : data_out = 24'b000000000000110111101100;
    16'b1111110010101101 : data_out = 24'b000000000000110111110000;
    16'b1111110010101110 : data_out = 24'b000000000000110111110011;
    16'b1111110010101111 : data_out = 24'b000000000000110111110111;
    16'b1111110010110000 : data_out = 24'b000000000000110111111010;
    16'b1111110010110001 : data_out = 24'b000000000000110111111110;
    16'b1111110010110010 : data_out = 24'b000000000000111000000001;
    16'b1111110010110011 : data_out = 24'b000000000000111000000101;
    16'b1111110010110100 : data_out = 24'b000000000000111000001000;
    16'b1111110010110101 : data_out = 24'b000000000000111000001100;
    16'b1111110010110110 : data_out = 24'b000000000000111000001111;
    16'b1111110010110111 : data_out = 24'b000000000000111000010011;
    16'b1111110010111000 : data_out = 24'b000000000000111000010110;
    16'b1111110010111001 : data_out = 24'b000000000000111000011010;
    16'b1111110010111010 : data_out = 24'b000000000000111000011101;
    16'b1111110010111011 : data_out = 24'b000000000000111000100001;
    16'b1111110010111100 : data_out = 24'b000000000000111000100101;
    16'b1111110010111101 : data_out = 24'b000000000000111000101000;
    16'b1111110010111110 : data_out = 24'b000000000000111000101100;
    16'b1111110010111111 : data_out = 24'b000000000000111000101111;
    16'b1111110011000000 : data_out = 24'b000000000000111000110011;
    16'b1111110011000001 : data_out = 24'b000000000000111000110110;
    16'b1111110011000010 : data_out = 24'b000000000000111000111010;
    16'b1111110011000011 : data_out = 24'b000000000000111000111101;
    16'b1111110011000100 : data_out = 24'b000000000000111001000001;
    16'b1111110011000101 : data_out = 24'b000000000000111001000100;
    16'b1111110011000110 : data_out = 24'b000000000000111001001000;
    16'b1111110011000111 : data_out = 24'b000000000000111001001100;
    16'b1111110011001000 : data_out = 24'b000000000000111001001111;
    16'b1111110011001001 : data_out = 24'b000000000000111001010011;
    16'b1111110011001010 : data_out = 24'b000000000000111001010110;
    16'b1111110011001011 : data_out = 24'b000000000000111001011010;
    16'b1111110011001100 : data_out = 24'b000000000000111001011110;
    16'b1111110011001101 : data_out = 24'b000000000000111001100001;
    16'b1111110011001110 : data_out = 24'b000000000000111001100101;
    16'b1111110011001111 : data_out = 24'b000000000000111001101000;
    16'b1111110011010000 : data_out = 24'b000000000000111001101100;
    16'b1111110011010001 : data_out = 24'b000000000000111001110000;
    16'b1111110011010010 : data_out = 24'b000000000000111001110011;
    16'b1111110011010011 : data_out = 24'b000000000000111001110111;
    16'b1111110011010100 : data_out = 24'b000000000000111001111010;
    16'b1111110011010101 : data_out = 24'b000000000000111001111110;
    16'b1111110011010110 : data_out = 24'b000000000000111010000010;
    16'b1111110011010111 : data_out = 24'b000000000000111010000101;
    16'b1111110011011000 : data_out = 24'b000000000000111010001001;
    16'b1111110011011001 : data_out = 24'b000000000000111010001101;
    16'b1111110011011010 : data_out = 24'b000000000000111010010000;
    16'b1111110011011011 : data_out = 24'b000000000000111010010100;
    16'b1111110011011100 : data_out = 24'b000000000000111010010111;
    16'b1111110011011101 : data_out = 24'b000000000000111010011011;
    16'b1111110011011110 : data_out = 24'b000000000000111010011111;
    16'b1111110011011111 : data_out = 24'b000000000000111010100010;
    16'b1111110011100000 : data_out = 24'b000000000000111010100110;
    16'b1111110011100001 : data_out = 24'b000000000000111010101010;
    16'b1111110011100010 : data_out = 24'b000000000000111010101101;
    16'b1111110011100011 : data_out = 24'b000000000000111010110001;
    16'b1111110011100100 : data_out = 24'b000000000000111010110101;
    16'b1111110011100101 : data_out = 24'b000000000000111010111000;
    16'b1111110011100110 : data_out = 24'b000000000000111010111100;
    16'b1111110011100111 : data_out = 24'b000000000000111011000000;
    16'b1111110011101000 : data_out = 24'b000000000000111011000011;
    16'b1111110011101001 : data_out = 24'b000000000000111011000111;
    16'b1111110011101010 : data_out = 24'b000000000000111011001011;
    16'b1111110011101011 : data_out = 24'b000000000000111011001111;
    16'b1111110011101100 : data_out = 24'b000000000000111011010010;
    16'b1111110011101101 : data_out = 24'b000000000000111011010110;
    16'b1111110011101110 : data_out = 24'b000000000000111011011010;
    16'b1111110011101111 : data_out = 24'b000000000000111011011101;
    16'b1111110011110000 : data_out = 24'b000000000000111011100001;
    16'b1111110011110001 : data_out = 24'b000000000000111011100101;
    16'b1111110011110010 : data_out = 24'b000000000000111011101001;
    16'b1111110011110011 : data_out = 24'b000000000000111011101100;
    16'b1111110011110100 : data_out = 24'b000000000000111011110000;
    16'b1111110011110101 : data_out = 24'b000000000000111011110100;
    16'b1111110011110110 : data_out = 24'b000000000000111011111000;
    16'b1111110011110111 : data_out = 24'b000000000000111011111011;
    16'b1111110011111000 : data_out = 24'b000000000000111011111111;
    16'b1111110011111001 : data_out = 24'b000000000000111100000011;
    16'b1111110011111010 : data_out = 24'b000000000000111100000111;
    16'b1111110011111011 : data_out = 24'b000000000000111100001010;
    16'b1111110011111100 : data_out = 24'b000000000000111100001110;
    16'b1111110011111101 : data_out = 24'b000000000000111100010010;
    16'b1111110011111110 : data_out = 24'b000000000000111100010110;
    16'b1111110011111111 : data_out = 24'b000000000000111100011001;
    16'b1111110100000000 : data_out = 24'b000000000000111100011101;
    16'b1111110100000001 : data_out = 24'b000000000000111100100001;
    16'b1111110100000010 : data_out = 24'b000000000000111100100101;
    16'b1111110100000011 : data_out = 24'b000000000000111100101000;
    16'b1111110100000100 : data_out = 24'b000000000000111100101100;
    16'b1111110100000101 : data_out = 24'b000000000000111100110000;
    16'b1111110100000110 : data_out = 24'b000000000000111100110100;
    16'b1111110100000111 : data_out = 24'b000000000000111100111000;
    16'b1111110100001000 : data_out = 24'b000000000000111100111011;
    16'b1111110100001001 : data_out = 24'b000000000000111100111111;
    16'b1111110100001010 : data_out = 24'b000000000000111101000011;
    16'b1111110100001011 : data_out = 24'b000000000000111101000111;
    16'b1111110100001100 : data_out = 24'b000000000000111101001011;
    16'b1111110100001101 : data_out = 24'b000000000000111101001111;
    16'b1111110100001110 : data_out = 24'b000000000000111101010010;
    16'b1111110100001111 : data_out = 24'b000000000000111101010110;
    16'b1111110100010000 : data_out = 24'b000000000000111101011010;
    16'b1111110100010001 : data_out = 24'b000000000000111101011110;
    16'b1111110100010010 : data_out = 24'b000000000000111101100010;
    16'b1111110100010011 : data_out = 24'b000000000000111101100110;
    16'b1111110100010100 : data_out = 24'b000000000000111101101001;
    16'b1111110100010101 : data_out = 24'b000000000000111101101101;
    16'b1111110100010110 : data_out = 24'b000000000000111101110001;
    16'b1111110100010111 : data_out = 24'b000000000000111101110101;
    16'b1111110100011000 : data_out = 24'b000000000000111101111001;
    16'b1111110100011001 : data_out = 24'b000000000000111101111101;
    16'b1111110100011010 : data_out = 24'b000000000000111110000001;
    16'b1111110100011011 : data_out = 24'b000000000000111110000101;
    16'b1111110100011100 : data_out = 24'b000000000000111110001000;
    16'b1111110100011101 : data_out = 24'b000000000000111110001100;
    16'b1111110100011110 : data_out = 24'b000000000000111110010000;
    16'b1111110100011111 : data_out = 24'b000000000000111110010100;
    16'b1111110100100000 : data_out = 24'b000000000000111110011000;
    16'b1111110100100001 : data_out = 24'b000000000000111110011100;
    16'b1111110100100010 : data_out = 24'b000000000000111110100000;
    16'b1111110100100011 : data_out = 24'b000000000000111110100100;
    16'b1111110100100100 : data_out = 24'b000000000000111110101000;
    16'b1111110100100101 : data_out = 24'b000000000000111110101100;
    16'b1111110100100110 : data_out = 24'b000000000000111110101111;
    16'b1111110100100111 : data_out = 24'b000000000000111110110011;
    16'b1111110100101000 : data_out = 24'b000000000000111110110111;
    16'b1111110100101001 : data_out = 24'b000000000000111110111011;
    16'b1111110100101010 : data_out = 24'b000000000000111110111111;
    16'b1111110100101011 : data_out = 24'b000000000000111111000011;
    16'b1111110100101100 : data_out = 24'b000000000000111111000111;
    16'b1111110100101101 : data_out = 24'b000000000000111111001011;
    16'b1111110100101110 : data_out = 24'b000000000000111111001111;
    16'b1111110100101111 : data_out = 24'b000000000000111111010011;
    16'b1111110100110000 : data_out = 24'b000000000000111111010111;
    16'b1111110100110001 : data_out = 24'b000000000000111111011011;
    16'b1111110100110010 : data_out = 24'b000000000000111111011111;
    16'b1111110100110011 : data_out = 24'b000000000000111111100011;
    16'b1111110100110100 : data_out = 24'b000000000000111111100111;
    16'b1111110100110101 : data_out = 24'b000000000000111111101011;
    16'b1111110100110110 : data_out = 24'b000000000000111111101111;
    16'b1111110100110111 : data_out = 24'b000000000000111111110011;
    16'b1111110100111000 : data_out = 24'b000000000000111111110111;
    16'b1111110100111001 : data_out = 24'b000000000000111111111011;
    16'b1111110100111010 : data_out = 24'b000000000000111111111111;
    16'b1111110100111011 : data_out = 24'b000000000001000000000011;
    16'b1111110100111100 : data_out = 24'b000000000001000000000111;
    16'b1111110100111101 : data_out = 24'b000000000001000000001011;
    16'b1111110100111110 : data_out = 24'b000000000001000000001111;
    16'b1111110100111111 : data_out = 24'b000000000001000000010011;
    16'b1111110101000000 : data_out = 24'b000000000001000000010111;
    16'b1111110101000001 : data_out = 24'b000000000001000000011011;
    16'b1111110101000010 : data_out = 24'b000000000001000000011111;
    16'b1111110101000011 : data_out = 24'b000000000001000000100011;
    16'b1111110101000100 : data_out = 24'b000000000001000000100111;
    16'b1111110101000101 : data_out = 24'b000000000001000000101011;
    16'b1111110101000110 : data_out = 24'b000000000001000000101111;
    16'b1111110101000111 : data_out = 24'b000000000001000000110011;
    16'b1111110101001000 : data_out = 24'b000000000001000000110111;
    16'b1111110101001001 : data_out = 24'b000000000001000000111011;
    16'b1111110101001010 : data_out = 24'b000000000001000000111111;
    16'b1111110101001011 : data_out = 24'b000000000001000001000011;
    16'b1111110101001100 : data_out = 24'b000000000001000001000111;
    16'b1111110101001101 : data_out = 24'b000000000001000001001011;
    16'b1111110101001110 : data_out = 24'b000000000001000001001111;
    16'b1111110101001111 : data_out = 24'b000000000001000001010011;
    16'b1111110101010000 : data_out = 24'b000000000001000001011000;
    16'b1111110101010001 : data_out = 24'b000000000001000001011100;
    16'b1111110101010010 : data_out = 24'b000000000001000001100000;
    16'b1111110101010011 : data_out = 24'b000000000001000001100100;
    16'b1111110101010100 : data_out = 24'b000000000001000001101000;
    16'b1111110101010101 : data_out = 24'b000000000001000001101100;
    16'b1111110101010110 : data_out = 24'b000000000001000001110000;
    16'b1111110101010111 : data_out = 24'b000000000001000001110100;
    16'b1111110101011000 : data_out = 24'b000000000001000001111000;
    16'b1111110101011001 : data_out = 24'b000000000001000001111101;
    16'b1111110101011010 : data_out = 24'b000000000001000010000001;
    16'b1111110101011011 : data_out = 24'b000000000001000010000101;
    16'b1111110101011100 : data_out = 24'b000000000001000010001001;
    16'b1111110101011101 : data_out = 24'b000000000001000010001101;
    16'b1111110101011110 : data_out = 24'b000000000001000010010001;
    16'b1111110101011111 : data_out = 24'b000000000001000010010101;
    16'b1111110101100000 : data_out = 24'b000000000001000010011001;
    16'b1111110101100001 : data_out = 24'b000000000001000010011110;
    16'b1111110101100010 : data_out = 24'b000000000001000010100010;
    16'b1111110101100011 : data_out = 24'b000000000001000010100110;
    16'b1111110101100100 : data_out = 24'b000000000001000010101010;
    16'b1111110101100101 : data_out = 24'b000000000001000010101110;
    16'b1111110101100110 : data_out = 24'b000000000001000010110010;
    16'b1111110101100111 : data_out = 24'b000000000001000010110111;
    16'b1111110101101000 : data_out = 24'b000000000001000010111011;
    16'b1111110101101001 : data_out = 24'b000000000001000010111111;
    16'b1111110101101010 : data_out = 24'b000000000001000011000011;
    16'b1111110101101011 : data_out = 24'b000000000001000011000111;
    16'b1111110101101100 : data_out = 24'b000000000001000011001100;
    16'b1111110101101101 : data_out = 24'b000000000001000011010000;
    16'b1111110101101110 : data_out = 24'b000000000001000011010100;
    16'b1111110101101111 : data_out = 24'b000000000001000011011000;
    16'b1111110101110000 : data_out = 24'b000000000001000011011100;
    16'b1111110101110001 : data_out = 24'b000000000001000011100001;
    16'b1111110101110010 : data_out = 24'b000000000001000011100101;
    16'b1111110101110011 : data_out = 24'b000000000001000011101001;
    16'b1111110101110100 : data_out = 24'b000000000001000011101101;
    16'b1111110101110101 : data_out = 24'b000000000001000011110010;
    16'b1111110101110110 : data_out = 24'b000000000001000011110110;
    16'b1111110101110111 : data_out = 24'b000000000001000011111010;
    16'b1111110101111000 : data_out = 24'b000000000001000011111110;
    16'b1111110101111001 : data_out = 24'b000000000001000100000010;
    16'b1111110101111010 : data_out = 24'b000000000001000100000111;
    16'b1111110101111011 : data_out = 24'b000000000001000100001011;
    16'b1111110101111100 : data_out = 24'b000000000001000100001111;
    16'b1111110101111101 : data_out = 24'b000000000001000100010100;
    16'b1111110101111110 : data_out = 24'b000000000001000100011000;
    16'b1111110101111111 : data_out = 24'b000000000001000100011100;
    16'b1111110110000000 : data_out = 24'b000000000001000100100000;
    16'b1111110110000001 : data_out = 24'b000000000001000100100101;
    16'b1111110110000010 : data_out = 24'b000000000001000100101001;
    16'b1111110110000011 : data_out = 24'b000000000001000100101101;
    16'b1111110110000100 : data_out = 24'b000000000001000100110010;
    16'b1111110110000101 : data_out = 24'b000000000001000100110110;
    16'b1111110110000110 : data_out = 24'b000000000001000100111010;
    16'b1111110110000111 : data_out = 24'b000000000001000100111110;
    16'b1111110110001000 : data_out = 24'b000000000001000101000011;
    16'b1111110110001001 : data_out = 24'b000000000001000101000111;
    16'b1111110110001010 : data_out = 24'b000000000001000101001011;
    16'b1111110110001011 : data_out = 24'b000000000001000101010000;
    16'b1111110110001100 : data_out = 24'b000000000001000101010100;
    16'b1111110110001101 : data_out = 24'b000000000001000101011000;
    16'b1111110110001110 : data_out = 24'b000000000001000101011101;
    16'b1111110110001111 : data_out = 24'b000000000001000101100001;
    16'b1111110110010000 : data_out = 24'b000000000001000101100101;
    16'b1111110110010001 : data_out = 24'b000000000001000101101010;
    16'b1111110110010010 : data_out = 24'b000000000001000101101110;
    16'b1111110110010011 : data_out = 24'b000000000001000101110010;
    16'b1111110110010100 : data_out = 24'b000000000001000101110111;
    16'b1111110110010101 : data_out = 24'b000000000001000101111011;
    16'b1111110110010110 : data_out = 24'b000000000001000110000000;
    16'b1111110110010111 : data_out = 24'b000000000001000110000100;
    16'b1111110110011000 : data_out = 24'b000000000001000110001000;
    16'b1111110110011001 : data_out = 24'b000000000001000110001101;
    16'b1111110110011010 : data_out = 24'b000000000001000110010001;
    16'b1111110110011011 : data_out = 24'b000000000001000110010110;
    16'b1111110110011100 : data_out = 24'b000000000001000110011010;
    16'b1111110110011101 : data_out = 24'b000000000001000110011110;
    16'b1111110110011110 : data_out = 24'b000000000001000110100011;
    16'b1111110110011111 : data_out = 24'b000000000001000110100111;
    16'b1111110110100000 : data_out = 24'b000000000001000110101100;
    16'b1111110110100001 : data_out = 24'b000000000001000110110000;
    16'b1111110110100010 : data_out = 24'b000000000001000110110100;
    16'b1111110110100011 : data_out = 24'b000000000001000110111001;
    16'b1111110110100100 : data_out = 24'b000000000001000110111101;
    16'b1111110110100101 : data_out = 24'b000000000001000111000010;
    16'b1111110110100110 : data_out = 24'b000000000001000111000110;
    16'b1111110110100111 : data_out = 24'b000000000001000111001011;
    16'b1111110110101000 : data_out = 24'b000000000001000111001111;
    16'b1111110110101001 : data_out = 24'b000000000001000111010011;
    16'b1111110110101010 : data_out = 24'b000000000001000111011000;
    16'b1111110110101011 : data_out = 24'b000000000001000111011100;
    16'b1111110110101100 : data_out = 24'b000000000001000111100001;
    16'b1111110110101101 : data_out = 24'b000000000001000111100101;
    16'b1111110110101110 : data_out = 24'b000000000001000111101010;
    16'b1111110110101111 : data_out = 24'b000000000001000111101110;
    16'b1111110110110000 : data_out = 24'b000000000001000111110011;
    16'b1111110110110001 : data_out = 24'b000000000001000111110111;
    16'b1111110110110010 : data_out = 24'b000000000001000111111100;
    16'b1111110110110011 : data_out = 24'b000000000001001000000000;
    16'b1111110110110100 : data_out = 24'b000000000001001000000101;
    16'b1111110110110101 : data_out = 24'b000000000001001000001001;
    16'b1111110110110110 : data_out = 24'b000000000001001000001110;
    16'b1111110110110111 : data_out = 24'b000000000001001000010010;
    16'b1111110110111000 : data_out = 24'b000000000001001000010111;
    16'b1111110110111001 : data_out = 24'b000000000001001000011011;
    16'b1111110110111010 : data_out = 24'b000000000001001000100000;
    16'b1111110110111011 : data_out = 24'b000000000001001000100100;
    16'b1111110110111100 : data_out = 24'b000000000001001000101001;
    16'b1111110110111101 : data_out = 24'b000000000001001000101110;
    16'b1111110110111110 : data_out = 24'b000000000001001000110010;
    16'b1111110110111111 : data_out = 24'b000000000001001000110111;
    16'b1111110111000000 : data_out = 24'b000000000001001000111011;
    16'b1111110111000001 : data_out = 24'b000000000001001001000000;
    16'b1111110111000010 : data_out = 24'b000000000001001001000100;
    16'b1111110111000011 : data_out = 24'b000000000001001001001001;
    16'b1111110111000100 : data_out = 24'b000000000001001001001101;
    16'b1111110111000101 : data_out = 24'b000000000001001001010010;
    16'b1111110111000110 : data_out = 24'b000000000001001001010111;
    16'b1111110111000111 : data_out = 24'b000000000001001001011011;
    16'b1111110111001000 : data_out = 24'b000000000001001001100000;
    16'b1111110111001001 : data_out = 24'b000000000001001001100100;
    16'b1111110111001010 : data_out = 24'b000000000001001001101001;
    16'b1111110111001011 : data_out = 24'b000000000001001001101110;
    16'b1111110111001100 : data_out = 24'b000000000001001001110010;
    16'b1111110111001101 : data_out = 24'b000000000001001001110111;
    16'b1111110111001110 : data_out = 24'b000000000001001001111011;
    16'b1111110111001111 : data_out = 24'b000000000001001010000000;
    16'b1111110111010000 : data_out = 24'b000000000001001010000101;
    16'b1111110111010001 : data_out = 24'b000000000001001010001001;
    16'b1111110111010010 : data_out = 24'b000000000001001010001110;
    16'b1111110111010011 : data_out = 24'b000000000001001010010011;
    16'b1111110111010100 : data_out = 24'b000000000001001010010111;
    16'b1111110111010101 : data_out = 24'b000000000001001010011100;
    16'b1111110111010110 : data_out = 24'b000000000001001010100001;
    16'b1111110111010111 : data_out = 24'b000000000001001010100101;
    16'b1111110111011000 : data_out = 24'b000000000001001010101010;
    16'b1111110111011001 : data_out = 24'b000000000001001010101111;
    16'b1111110111011010 : data_out = 24'b000000000001001010110011;
    16'b1111110111011011 : data_out = 24'b000000000001001010111000;
    16'b1111110111011100 : data_out = 24'b000000000001001010111101;
    16'b1111110111011101 : data_out = 24'b000000000001001011000001;
    16'b1111110111011110 : data_out = 24'b000000000001001011000110;
    16'b1111110111011111 : data_out = 24'b000000000001001011001011;
    16'b1111110111100000 : data_out = 24'b000000000001001011001111;
    16'b1111110111100001 : data_out = 24'b000000000001001011010100;
    16'b1111110111100010 : data_out = 24'b000000000001001011011001;
    16'b1111110111100011 : data_out = 24'b000000000001001011011101;
    16'b1111110111100100 : data_out = 24'b000000000001001011100010;
    16'b1111110111100101 : data_out = 24'b000000000001001011100111;
    16'b1111110111100110 : data_out = 24'b000000000001001011101100;
    16'b1111110111100111 : data_out = 24'b000000000001001011110000;
    16'b1111110111101000 : data_out = 24'b000000000001001011110101;
    16'b1111110111101001 : data_out = 24'b000000000001001011111010;
    16'b1111110111101010 : data_out = 24'b000000000001001011111111;
    16'b1111110111101011 : data_out = 24'b000000000001001100000011;
    16'b1111110111101100 : data_out = 24'b000000000001001100001000;
    16'b1111110111101101 : data_out = 24'b000000000001001100001101;
    16'b1111110111101110 : data_out = 24'b000000000001001100010010;
    16'b1111110111101111 : data_out = 24'b000000000001001100010110;
    16'b1111110111110000 : data_out = 24'b000000000001001100011011;
    16'b1111110111110001 : data_out = 24'b000000000001001100100000;
    16'b1111110111110010 : data_out = 24'b000000000001001100100101;
    16'b1111110111110011 : data_out = 24'b000000000001001100101010;
    16'b1111110111110100 : data_out = 24'b000000000001001100101110;
    16'b1111110111110101 : data_out = 24'b000000000001001100110011;
    16'b1111110111110110 : data_out = 24'b000000000001001100111000;
    16'b1111110111110111 : data_out = 24'b000000000001001100111101;
    16'b1111110111111000 : data_out = 24'b000000000001001101000010;
    16'b1111110111111001 : data_out = 24'b000000000001001101000110;
    16'b1111110111111010 : data_out = 24'b000000000001001101001011;
    16'b1111110111111011 : data_out = 24'b000000000001001101010000;
    16'b1111110111111100 : data_out = 24'b000000000001001101010101;
    16'b1111110111111101 : data_out = 24'b000000000001001101011010;
    16'b1111110111111110 : data_out = 24'b000000000001001101011111;
    16'b1111110111111111 : data_out = 24'b000000000001001101100011;
    16'b1111111000000000 : data_out = 24'b000000000001001101101000;
    16'b1111111000000001 : data_out = 24'b000000000001001101101101;
    16'b1111111000000010 : data_out = 24'b000000000001001101110010;
    16'b1111111000000011 : data_out = 24'b000000000001001101110111;
    16'b1111111000000100 : data_out = 24'b000000000001001101111100;
    16'b1111111000000101 : data_out = 24'b000000000001001110000001;
    16'b1111111000000110 : data_out = 24'b000000000001001110000101;
    16'b1111111000000111 : data_out = 24'b000000000001001110001010;
    16'b1111111000001000 : data_out = 24'b000000000001001110001111;
    16'b1111111000001001 : data_out = 24'b000000000001001110010100;
    16'b1111111000001010 : data_out = 24'b000000000001001110011001;
    16'b1111111000001011 : data_out = 24'b000000000001001110011110;
    16'b1111111000001100 : data_out = 24'b000000000001001110100011;
    16'b1111111000001101 : data_out = 24'b000000000001001110101000;
    16'b1111111000001110 : data_out = 24'b000000000001001110101101;
    16'b1111111000001111 : data_out = 24'b000000000001001110110010;
    16'b1111111000010000 : data_out = 24'b000000000001001110110110;
    16'b1111111000010001 : data_out = 24'b000000000001001110111011;
    16'b1111111000010010 : data_out = 24'b000000000001001111000000;
    16'b1111111000010011 : data_out = 24'b000000000001001111000101;
    16'b1111111000010100 : data_out = 24'b000000000001001111001010;
    16'b1111111000010101 : data_out = 24'b000000000001001111001111;
    16'b1111111000010110 : data_out = 24'b000000000001001111010100;
    16'b1111111000010111 : data_out = 24'b000000000001001111011001;
    16'b1111111000011000 : data_out = 24'b000000000001001111011110;
    16'b1111111000011001 : data_out = 24'b000000000001001111100011;
    16'b1111111000011010 : data_out = 24'b000000000001001111101000;
    16'b1111111000011011 : data_out = 24'b000000000001001111101101;
    16'b1111111000011100 : data_out = 24'b000000000001001111110010;
    16'b1111111000011101 : data_out = 24'b000000000001001111110111;
    16'b1111111000011110 : data_out = 24'b000000000001001111111100;
    16'b1111111000011111 : data_out = 24'b000000000001010000000001;
    16'b1111111000100000 : data_out = 24'b000000000001010000000110;
    16'b1111111000100001 : data_out = 24'b000000000001010000001011;
    16'b1111111000100010 : data_out = 24'b000000000001010000010000;
    16'b1111111000100011 : data_out = 24'b000000000001010000010101;
    16'b1111111000100100 : data_out = 24'b000000000001010000011010;
    16'b1111111000100101 : data_out = 24'b000000000001010000011111;
    16'b1111111000100110 : data_out = 24'b000000000001010000100100;
    16'b1111111000100111 : data_out = 24'b000000000001010000101001;
    16'b1111111000101000 : data_out = 24'b000000000001010000101110;
    16'b1111111000101001 : data_out = 24'b000000000001010000110011;
    16'b1111111000101010 : data_out = 24'b000000000001010000111000;
    16'b1111111000101011 : data_out = 24'b000000000001010000111101;
    16'b1111111000101100 : data_out = 24'b000000000001010001000010;
    16'b1111111000101101 : data_out = 24'b000000000001010001000111;
    16'b1111111000101110 : data_out = 24'b000000000001010001001100;
    16'b1111111000101111 : data_out = 24'b000000000001010001010010;
    16'b1111111000110000 : data_out = 24'b000000000001010001010111;
    16'b1111111000110001 : data_out = 24'b000000000001010001011100;
    16'b1111111000110010 : data_out = 24'b000000000001010001100001;
    16'b1111111000110011 : data_out = 24'b000000000001010001100110;
    16'b1111111000110100 : data_out = 24'b000000000001010001101011;
    16'b1111111000110101 : data_out = 24'b000000000001010001110000;
    16'b1111111000110110 : data_out = 24'b000000000001010001110101;
    16'b1111111000110111 : data_out = 24'b000000000001010001111010;
    16'b1111111000111000 : data_out = 24'b000000000001010001111111;
    16'b1111111000111001 : data_out = 24'b000000000001010010000101;
    16'b1111111000111010 : data_out = 24'b000000000001010010001010;
    16'b1111111000111011 : data_out = 24'b000000000001010010001111;
    16'b1111111000111100 : data_out = 24'b000000000001010010010100;
    16'b1111111000111101 : data_out = 24'b000000000001010010011001;
    16'b1111111000111110 : data_out = 24'b000000000001010010011110;
    16'b1111111000111111 : data_out = 24'b000000000001010010100011;
    16'b1111111001000000 : data_out = 24'b000000000001010010101001;
    16'b1111111001000001 : data_out = 24'b000000000001010010101110;
    16'b1111111001000010 : data_out = 24'b000000000001010010110011;
    16'b1111111001000011 : data_out = 24'b000000000001010010111000;
    16'b1111111001000100 : data_out = 24'b000000000001010010111101;
    16'b1111111001000101 : data_out = 24'b000000000001010011000011;
    16'b1111111001000110 : data_out = 24'b000000000001010011001000;
    16'b1111111001000111 : data_out = 24'b000000000001010011001101;
    16'b1111111001001000 : data_out = 24'b000000000001010011010010;
    16'b1111111001001001 : data_out = 24'b000000000001010011010111;
    16'b1111111001001010 : data_out = 24'b000000000001010011011101;
    16'b1111111001001011 : data_out = 24'b000000000001010011100010;
    16'b1111111001001100 : data_out = 24'b000000000001010011100111;
    16'b1111111001001101 : data_out = 24'b000000000001010011101100;
    16'b1111111001001110 : data_out = 24'b000000000001010011110001;
    16'b1111111001001111 : data_out = 24'b000000000001010011110111;
    16'b1111111001010000 : data_out = 24'b000000000001010011111100;
    16'b1111111001010001 : data_out = 24'b000000000001010100000001;
    16'b1111111001010010 : data_out = 24'b000000000001010100000110;
    16'b1111111001010011 : data_out = 24'b000000000001010100001100;
    16'b1111111001010100 : data_out = 24'b000000000001010100010001;
    16'b1111111001010101 : data_out = 24'b000000000001010100010110;
    16'b1111111001010110 : data_out = 24'b000000000001010100011100;
    16'b1111111001010111 : data_out = 24'b000000000001010100100001;
    16'b1111111001011000 : data_out = 24'b000000000001010100100110;
    16'b1111111001011001 : data_out = 24'b000000000001010100101011;
    16'b1111111001011010 : data_out = 24'b000000000001010100110001;
    16'b1111111001011011 : data_out = 24'b000000000001010100110110;
    16'b1111111001011100 : data_out = 24'b000000000001010100111011;
    16'b1111111001011101 : data_out = 24'b000000000001010101000001;
    16'b1111111001011110 : data_out = 24'b000000000001010101000110;
    16'b1111111001011111 : data_out = 24'b000000000001010101001011;
    16'b1111111001100000 : data_out = 24'b000000000001010101010001;
    16'b1111111001100001 : data_out = 24'b000000000001010101010110;
    16'b1111111001100010 : data_out = 24'b000000000001010101011011;
    16'b1111111001100011 : data_out = 24'b000000000001010101100001;
    16'b1111111001100100 : data_out = 24'b000000000001010101100110;
    16'b1111111001100101 : data_out = 24'b000000000001010101101011;
    16'b1111111001100110 : data_out = 24'b000000000001010101110001;
    16'b1111111001100111 : data_out = 24'b000000000001010101110110;
    16'b1111111001101000 : data_out = 24'b000000000001010101111011;
    16'b1111111001101001 : data_out = 24'b000000000001010110000001;
    16'b1111111001101010 : data_out = 24'b000000000001010110000110;
    16'b1111111001101011 : data_out = 24'b000000000001010110001011;
    16'b1111111001101100 : data_out = 24'b000000000001010110010001;
    16'b1111111001101101 : data_out = 24'b000000000001010110010110;
    16'b1111111001101110 : data_out = 24'b000000000001010110011100;
    16'b1111111001101111 : data_out = 24'b000000000001010110100001;
    16'b1111111001110000 : data_out = 24'b000000000001010110100110;
    16'b1111111001110001 : data_out = 24'b000000000001010110101100;
    16'b1111111001110010 : data_out = 24'b000000000001010110110001;
    16'b1111111001110011 : data_out = 24'b000000000001010110110111;
    16'b1111111001110100 : data_out = 24'b000000000001010110111100;
    16'b1111111001110101 : data_out = 24'b000000000001010111000010;
    16'b1111111001110110 : data_out = 24'b000000000001010111000111;
    16'b1111111001110111 : data_out = 24'b000000000001010111001101;
    16'b1111111001111000 : data_out = 24'b000000000001010111010010;
    16'b1111111001111001 : data_out = 24'b000000000001010111010111;
    16'b1111111001111010 : data_out = 24'b000000000001010111011101;
    16'b1111111001111011 : data_out = 24'b000000000001010111100010;
    16'b1111111001111100 : data_out = 24'b000000000001010111101000;
    16'b1111111001111101 : data_out = 24'b000000000001010111101101;
    16'b1111111001111110 : data_out = 24'b000000000001010111110011;
    16'b1111111001111111 : data_out = 24'b000000000001010111111000;
    16'b1111111010000000 : data_out = 24'b000000000001010111111110;
    16'b1111111010000001 : data_out = 24'b000000000001011000000011;
    16'b1111111010000010 : data_out = 24'b000000000001011000001001;
    16'b1111111010000011 : data_out = 24'b000000000001011000001110;
    16'b1111111010000100 : data_out = 24'b000000000001011000010100;
    16'b1111111010000101 : data_out = 24'b000000000001011000011001;
    16'b1111111010000110 : data_out = 24'b000000000001011000011111;
    16'b1111111010000111 : data_out = 24'b000000000001011000100100;
    16'b1111111010001000 : data_out = 24'b000000000001011000101010;
    16'b1111111010001001 : data_out = 24'b000000000001011000101111;
    16'b1111111010001010 : data_out = 24'b000000000001011000110101;
    16'b1111111010001011 : data_out = 24'b000000000001011000111011;
    16'b1111111010001100 : data_out = 24'b000000000001011001000000;
    16'b1111111010001101 : data_out = 24'b000000000001011001000110;
    16'b1111111010001110 : data_out = 24'b000000000001011001001011;
    16'b1111111010001111 : data_out = 24'b000000000001011001010001;
    16'b1111111010010000 : data_out = 24'b000000000001011001010110;
    16'b1111111010010001 : data_out = 24'b000000000001011001011100;
    16'b1111111010010010 : data_out = 24'b000000000001011001100010;
    16'b1111111010010011 : data_out = 24'b000000000001011001100111;
    16'b1111111010010100 : data_out = 24'b000000000001011001101101;
    16'b1111111010010101 : data_out = 24'b000000000001011001110010;
    16'b1111111010010110 : data_out = 24'b000000000001011001111000;
    16'b1111111010010111 : data_out = 24'b000000000001011001111110;
    16'b1111111010011000 : data_out = 24'b000000000001011010000011;
    16'b1111111010011001 : data_out = 24'b000000000001011010001001;
    16'b1111111010011010 : data_out = 24'b000000000001011010001111;
    16'b1111111010011011 : data_out = 24'b000000000001011010010100;
    16'b1111111010011100 : data_out = 24'b000000000001011010011010;
    16'b1111111010011101 : data_out = 24'b000000000001011010100000;
    16'b1111111010011110 : data_out = 24'b000000000001011010100101;
    16'b1111111010011111 : data_out = 24'b000000000001011010101011;
    16'b1111111010100000 : data_out = 24'b000000000001011010110000;
    16'b1111111010100001 : data_out = 24'b000000000001011010110110;
    16'b1111111010100010 : data_out = 24'b000000000001011010111100;
    16'b1111111010100011 : data_out = 24'b000000000001011011000010;
    16'b1111111010100100 : data_out = 24'b000000000001011011000111;
    16'b1111111010100101 : data_out = 24'b000000000001011011001101;
    16'b1111111010100110 : data_out = 24'b000000000001011011010011;
    16'b1111111010100111 : data_out = 24'b000000000001011011011000;
    16'b1111111010101000 : data_out = 24'b000000000001011011011110;
    16'b1111111010101001 : data_out = 24'b000000000001011011100100;
    16'b1111111010101010 : data_out = 24'b000000000001011011101010;
    16'b1111111010101011 : data_out = 24'b000000000001011011101111;
    16'b1111111010101100 : data_out = 24'b000000000001011011110101;
    16'b1111111010101101 : data_out = 24'b000000000001011011111011;
    16'b1111111010101110 : data_out = 24'b000000000001011100000000;
    16'b1111111010101111 : data_out = 24'b000000000001011100000110;
    16'b1111111010110000 : data_out = 24'b000000000001011100001100;
    16'b1111111010110001 : data_out = 24'b000000000001011100010010;
    16'b1111111010110010 : data_out = 24'b000000000001011100011000;
    16'b1111111010110011 : data_out = 24'b000000000001011100011101;
    16'b1111111010110100 : data_out = 24'b000000000001011100100011;
    16'b1111111010110101 : data_out = 24'b000000000001011100101001;
    16'b1111111010110110 : data_out = 24'b000000000001011100101111;
    16'b1111111010110111 : data_out = 24'b000000000001011100110100;
    16'b1111111010111000 : data_out = 24'b000000000001011100111010;
    16'b1111111010111001 : data_out = 24'b000000000001011101000000;
    16'b1111111010111010 : data_out = 24'b000000000001011101000110;
    16'b1111111010111011 : data_out = 24'b000000000001011101001100;
    16'b1111111010111100 : data_out = 24'b000000000001011101010010;
    16'b1111111010111101 : data_out = 24'b000000000001011101010111;
    16'b1111111010111110 : data_out = 24'b000000000001011101011101;
    16'b1111111010111111 : data_out = 24'b000000000001011101100011;
    16'b1111111011000000 : data_out = 24'b000000000001011101101001;
    16'b1111111011000001 : data_out = 24'b000000000001011101101111;
    16'b1111111011000010 : data_out = 24'b000000000001011101110101;
    16'b1111111011000011 : data_out = 24'b000000000001011101111010;
    16'b1111111011000100 : data_out = 24'b000000000001011110000000;
    16'b1111111011000101 : data_out = 24'b000000000001011110000110;
    16'b1111111011000110 : data_out = 24'b000000000001011110001100;
    16'b1111111011000111 : data_out = 24'b000000000001011110010010;
    16'b1111111011001000 : data_out = 24'b000000000001011110011000;
    16'b1111111011001001 : data_out = 24'b000000000001011110011110;
    16'b1111111011001010 : data_out = 24'b000000000001011110100100;
    16'b1111111011001011 : data_out = 24'b000000000001011110101010;
    16'b1111111011001100 : data_out = 24'b000000000001011110110000;
    16'b1111111011001101 : data_out = 24'b000000000001011110110101;
    16'b1111111011001110 : data_out = 24'b000000000001011110111011;
    16'b1111111011001111 : data_out = 24'b000000000001011111000001;
    16'b1111111011010000 : data_out = 24'b000000000001011111000111;
    16'b1111111011010001 : data_out = 24'b000000000001011111001101;
    16'b1111111011010010 : data_out = 24'b000000000001011111010011;
    16'b1111111011010011 : data_out = 24'b000000000001011111011001;
    16'b1111111011010100 : data_out = 24'b000000000001011111011111;
    16'b1111111011010101 : data_out = 24'b000000000001011111100101;
    16'b1111111011010110 : data_out = 24'b000000000001011111101011;
    16'b1111111011010111 : data_out = 24'b000000000001011111110001;
    16'b1111111011011000 : data_out = 24'b000000000001011111110111;
    16'b1111111011011001 : data_out = 24'b000000000001011111111101;
    16'b1111111011011010 : data_out = 24'b000000000001100000000011;
    16'b1111111011011011 : data_out = 24'b000000000001100000001001;
    16'b1111111011011100 : data_out = 24'b000000000001100000001111;
    16'b1111111011011101 : data_out = 24'b000000000001100000010101;
    16'b1111111011011110 : data_out = 24'b000000000001100000011011;
    16'b1111111011011111 : data_out = 24'b000000000001100000100001;
    16'b1111111011100000 : data_out = 24'b000000000001100000100111;
    16'b1111111011100001 : data_out = 24'b000000000001100000101101;
    16'b1111111011100010 : data_out = 24'b000000000001100000110011;
    16'b1111111011100011 : data_out = 24'b000000000001100000111001;
    16'b1111111011100100 : data_out = 24'b000000000001100000111111;
    16'b1111111011100101 : data_out = 24'b000000000001100001000101;
    16'b1111111011100110 : data_out = 24'b000000000001100001001011;
    16'b1111111011100111 : data_out = 24'b000000000001100001010010;
    16'b1111111011101000 : data_out = 24'b000000000001100001011000;
    16'b1111111011101001 : data_out = 24'b000000000001100001011110;
    16'b1111111011101010 : data_out = 24'b000000000001100001100100;
    16'b1111111011101011 : data_out = 24'b000000000001100001101010;
    16'b1111111011101100 : data_out = 24'b000000000001100001110000;
    16'b1111111011101101 : data_out = 24'b000000000001100001110110;
    16'b1111111011101110 : data_out = 24'b000000000001100001111100;
    16'b1111111011101111 : data_out = 24'b000000000001100010000010;
    16'b1111111011110000 : data_out = 24'b000000000001100010001001;
    16'b1111111011110001 : data_out = 24'b000000000001100010001111;
    16'b1111111011110010 : data_out = 24'b000000000001100010010101;
    16'b1111111011110011 : data_out = 24'b000000000001100010011011;
    16'b1111111011110100 : data_out = 24'b000000000001100010100001;
    16'b1111111011110101 : data_out = 24'b000000000001100010100111;
    16'b1111111011110110 : data_out = 24'b000000000001100010101101;
    16'b1111111011110111 : data_out = 24'b000000000001100010110100;
    16'b1111111011111000 : data_out = 24'b000000000001100010111010;
    16'b1111111011111001 : data_out = 24'b000000000001100011000000;
    16'b1111111011111010 : data_out = 24'b000000000001100011000110;
    16'b1111111011111011 : data_out = 24'b000000000001100011001100;
    16'b1111111011111100 : data_out = 24'b000000000001100011010011;
    16'b1111111011111101 : data_out = 24'b000000000001100011011001;
    16'b1111111011111110 : data_out = 24'b000000000001100011011111;
    16'b1111111011111111 : data_out = 24'b000000000001100011100101;
    16'b1111111100000000 : data_out = 24'b000000000001100011101011;
    16'b1111111100000001 : data_out = 24'b000000000001100011110010;
    16'b1111111100000010 : data_out = 24'b000000000001100011111000;
    16'b1111111100000011 : data_out = 24'b000000000001100011111110;
    16'b1111111100000100 : data_out = 24'b000000000001100100000100;
    16'b1111111100000101 : data_out = 24'b000000000001100100001011;
    16'b1111111100000110 : data_out = 24'b000000000001100100010001;
    16'b1111111100000111 : data_out = 24'b000000000001100100010111;
    16'b1111111100001000 : data_out = 24'b000000000001100100011101;
    16'b1111111100001001 : data_out = 24'b000000000001100100100100;
    16'b1111111100001010 : data_out = 24'b000000000001100100101010;
    16'b1111111100001011 : data_out = 24'b000000000001100100110000;
    16'b1111111100001100 : data_out = 24'b000000000001100100110111;
    16'b1111111100001101 : data_out = 24'b000000000001100100111101;
    16'b1111111100001110 : data_out = 24'b000000000001100101000011;
    16'b1111111100001111 : data_out = 24'b000000000001100101001010;
    16'b1111111100010000 : data_out = 24'b000000000001100101010000;
    16'b1111111100010001 : data_out = 24'b000000000001100101010110;
    16'b1111111100010010 : data_out = 24'b000000000001100101011101;
    16'b1111111100010011 : data_out = 24'b000000000001100101100011;
    16'b1111111100010100 : data_out = 24'b000000000001100101101001;
    16'b1111111100010101 : data_out = 24'b000000000001100101110000;
    16'b1111111100010110 : data_out = 24'b000000000001100101110110;
    16'b1111111100010111 : data_out = 24'b000000000001100101111100;
    16'b1111111100011000 : data_out = 24'b000000000001100110000011;
    16'b1111111100011001 : data_out = 24'b000000000001100110001001;
    16'b1111111100011010 : data_out = 24'b000000000001100110010000;
    16'b1111111100011011 : data_out = 24'b000000000001100110010110;
    16'b1111111100011100 : data_out = 24'b000000000001100110011100;
    16'b1111111100011101 : data_out = 24'b000000000001100110100011;
    16'b1111111100011110 : data_out = 24'b000000000001100110101001;
    16'b1111111100011111 : data_out = 24'b000000000001100110110000;
    16'b1111111100100000 : data_out = 24'b000000000001100110110110;
    16'b1111111100100001 : data_out = 24'b000000000001100110111100;
    16'b1111111100100010 : data_out = 24'b000000000001100111000011;
    16'b1111111100100011 : data_out = 24'b000000000001100111001001;
    16'b1111111100100100 : data_out = 24'b000000000001100111010000;
    16'b1111111100100101 : data_out = 24'b000000000001100111010110;
    16'b1111111100100110 : data_out = 24'b000000000001100111011101;
    16'b1111111100100111 : data_out = 24'b000000000001100111100011;
    16'b1111111100101000 : data_out = 24'b000000000001100111101010;
    16'b1111111100101001 : data_out = 24'b000000000001100111110000;
    16'b1111111100101010 : data_out = 24'b000000000001100111110111;
    16'b1111111100101011 : data_out = 24'b000000000001100111111101;
    16'b1111111100101100 : data_out = 24'b000000000001101000000100;
    16'b1111111100101101 : data_out = 24'b000000000001101000001010;
    16'b1111111100101110 : data_out = 24'b000000000001101000010001;
    16'b1111111100101111 : data_out = 24'b000000000001101000010111;
    16'b1111111100110000 : data_out = 24'b000000000001101000011110;
    16'b1111111100110001 : data_out = 24'b000000000001101000100100;
    16'b1111111100110010 : data_out = 24'b000000000001101000101011;
    16'b1111111100110011 : data_out = 24'b000000000001101000110001;
    16'b1111111100110100 : data_out = 24'b000000000001101000111000;
    16'b1111111100110101 : data_out = 24'b000000000001101000111110;
    16'b1111111100110110 : data_out = 24'b000000000001101001000101;
    16'b1111111100110111 : data_out = 24'b000000000001101001001011;
    16'b1111111100111000 : data_out = 24'b000000000001101001010010;
    16'b1111111100111001 : data_out = 24'b000000000001101001011001;
    16'b1111111100111010 : data_out = 24'b000000000001101001011111;
    16'b1111111100111011 : data_out = 24'b000000000001101001100110;
    16'b1111111100111100 : data_out = 24'b000000000001101001101100;
    16'b1111111100111101 : data_out = 24'b000000000001101001110011;
    16'b1111111100111110 : data_out = 24'b000000000001101001111010;
    16'b1111111100111111 : data_out = 24'b000000000001101010000000;
    16'b1111111101000000 : data_out = 24'b000000000001101010000111;
    16'b1111111101000001 : data_out = 24'b000000000001101010001110;
    16'b1111111101000010 : data_out = 24'b000000000001101010010100;
    16'b1111111101000011 : data_out = 24'b000000000001101010011011;
    16'b1111111101000100 : data_out = 24'b000000000001101010100001;
    16'b1111111101000101 : data_out = 24'b000000000001101010101000;
    16'b1111111101000110 : data_out = 24'b000000000001101010101111;
    16'b1111111101000111 : data_out = 24'b000000000001101010110101;
    16'b1111111101001000 : data_out = 24'b000000000001101010111100;
    16'b1111111101001001 : data_out = 24'b000000000001101011000011;
    16'b1111111101001010 : data_out = 24'b000000000001101011001010;
    16'b1111111101001011 : data_out = 24'b000000000001101011010000;
    16'b1111111101001100 : data_out = 24'b000000000001101011010111;
    16'b1111111101001101 : data_out = 24'b000000000001101011011110;
    16'b1111111101001110 : data_out = 24'b000000000001101011100100;
    16'b1111111101001111 : data_out = 24'b000000000001101011101011;
    16'b1111111101010000 : data_out = 24'b000000000001101011110010;
    16'b1111111101010001 : data_out = 24'b000000000001101011111001;
    16'b1111111101010010 : data_out = 24'b000000000001101011111111;
    16'b1111111101010011 : data_out = 24'b000000000001101100000110;
    16'b1111111101010100 : data_out = 24'b000000000001101100001101;
    16'b1111111101010101 : data_out = 24'b000000000001101100010100;
    16'b1111111101010110 : data_out = 24'b000000000001101100011010;
    16'b1111111101010111 : data_out = 24'b000000000001101100100001;
    16'b1111111101011000 : data_out = 24'b000000000001101100101000;
    16'b1111111101011001 : data_out = 24'b000000000001101100101111;
    16'b1111111101011010 : data_out = 24'b000000000001101100110110;
    16'b1111111101011011 : data_out = 24'b000000000001101100111100;
    16'b1111111101011100 : data_out = 24'b000000000001101101000011;
    16'b1111111101011101 : data_out = 24'b000000000001101101001010;
    16'b1111111101011110 : data_out = 24'b000000000001101101010001;
    16'b1111111101011111 : data_out = 24'b000000000001101101011000;
    16'b1111111101100000 : data_out = 24'b000000000001101101011110;
    16'b1111111101100001 : data_out = 24'b000000000001101101100101;
    16'b1111111101100010 : data_out = 24'b000000000001101101101100;
    16'b1111111101100011 : data_out = 24'b000000000001101101110011;
    16'b1111111101100100 : data_out = 24'b000000000001101101111010;
    16'b1111111101100101 : data_out = 24'b000000000001101110000001;
    16'b1111111101100110 : data_out = 24'b000000000001101110001000;
    16'b1111111101100111 : data_out = 24'b000000000001101110001111;
    16'b1111111101101000 : data_out = 24'b000000000001101110010101;
    16'b1111111101101001 : data_out = 24'b000000000001101110011100;
    16'b1111111101101010 : data_out = 24'b000000000001101110100011;
    16'b1111111101101011 : data_out = 24'b000000000001101110101010;
    16'b1111111101101100 : data_out = 24'b000000000001101110110001;
    16'b1111111101101101 : data_out = 24'b000000000001101110111000;
    16'b1111111101101110 : data_out = 24'b000000000001101110111111;
    16'b1111111101101111 : data_out = 24'b000000000001101111000110;
    16'b1111111101110000 : data_out = 24'b000000000001101111001101;
    16'b1111111101110001 : data_out = 24'b000000000001101111010100;
    16'b1111111101110010 : data_out = 24'b000000000001101111011011;
    16'b1111111101110011 : data_out = 24'b000000000001101111100010;
    16'b1111111101110100 : data_out = 24'b000000000001101111101001;
    16'b1111111101110101 : data_out = 24'b000000000001101111110000;
    16'b1111111101110110 : data_out = 24'b000000000001101111110111;
    16'b1111111101110111 : data_out = 24'b000000000001101111111110;
    16'b1111111101111000 : data_out = 24'b000000000001110000000101;
    16'b1111111101111001 : data_out = 24'b000000000001110000001100;
    16'b1111111101111010 : data_out = 24'b000000000001110000010011;
    16'b1111111101111011 : data_out = 24'b000000000001110000011010;
    16'b1111111101111100 : data_out = 24'b000000000001110000100001;
    16'b1111111101111101 : data_out = 24'b000000000001110000101000;
    16'b1111111101111110 : data_out = 24'b000000000001110000101111;
    16'b1111111101111111 : data_out = 24'b000000000001110000110110;
    16'b1111111110000000 : data_out = 24'b000000000001110000111101;
    16'b1111111110000001 : data_out = 24'b000000000001110001000100;
    16'b1111111110000010 : data_out = 24'b000000000001110001001011;
    16'b1111111110000011 : data_out = 24'b000000000001110001010010;
    16'b1111111110000100 : data_out = 24'b000000000001110001011001;
    16'b1111111110000101 : data_out = 24'b000000000001110001100000;
    16'b1111111110000110 : data_out = 24'b000000000001110001100111;
    16'b1111111110000111 : data_out = 24'b000000000001110001101111;
    16'b1111111110001000 : data_out = 24'b000000000001110001110110;
    16'b1111111110001001 : data_out = 24'b000000000001110001111101;
    16'b1111111110001010 : data_out = 24'b000000000001110010000100;
    16'b1111111110001011 : data_out = 24'b000000000001110010001011;
    16'b1111111110001100 : data_out = 24'b000000000001110010010010;
    16'b1111111110001101 : data_out = 24'b000000000001110010011001;
    16'b1111111110001110 : data_out = 24'b000000000001110010100000;
    16'b1111111110001111 : data_out = 24'b000000000001110010101000;
    16'b1111111110010000 : data_out = 24'b000000000001110010101111;
    16'b1111111110010001 : data_out = 24'b000000000001110010110110;
    16'b1111111110010010 : data_out = 24'b000000000001110010111101;
    16'b1111111110010011 : data_out = 24'b000000000001110011000100;
    16'b1111111110010100 : data_out = 24'b000000000001110011001100;
    16'b1111111110010101 : data_out = 24'b000000000001110011010011;
    16'b1111111110010110 : data_out = 24'b000000000001110011011010;
    16'b1111111110010111 : data_out = 24'b000000000001110011100001;
    16'b1111111110011000 : data_out = 24'b000000000001110011101000;
    16'b1111111110011001 : data_out = 24'b000000000001110011110000;
    16'b1111111110011010 : data_out = 24'b000000000001110011110111;
    16'b1111111110011011 : data_out = 24'b000000000001110011111110;
    16'b1111111110011100 : data_out = 24'b000000000001110100000101;
    16'b1111111110011101 : data_out = 24'b000000000001110100001101;
    16'b1111111110011110 : data_out = 24'b000000000001110100010100;
    16'b1111111110011111 : data_out = 24'b000000000001110100011011;
    16'b1111111110100000 : data_out = 24'b000000000001110100100010;
    16'b1111111110100001 : data_out = 24'b000000000001110100101010;
    16'b1111111110100010 : data_out = 24'b000000000001110100110001;
    16'b1111111110100011 : data_out = 24'b000000000001110100111000;
    16'b1111111110100100 : data_out = 24'b000000000001110101000000;
    16'b1111111110100101 : data_out = 24'b000000000001110101000111;
    16'b1111111110100110 : data_out = 24'b000000000001110101001110;
    16'b1111111110100111 : data_out = 24'b000000000001110101010110;
    16'b1111111110101000 : data_out = 24'b000000000001110101011101;
    16'b1111111110101001 : data_out = 24'b000000000001110101100100;
    16'b1111111110101010 : data_out = 24'b000000000001110101101100;
    16'b1111111110101011 : data_out = 24'b000000000001110101110011;
    16'b1111111110101100 : data_out = 24'b000000000001110101111010;
    16'b1111111110101101 : data_out = 24'b000000000001110110000010;
    16'b1111111110101110 : data_out = 24'b000000000001110110001001;
    16'b1111111110101111 : data_out = 24'b000000000001110110010000;
    16'b1111111110110000 : data_out = 24'b000000000001110110011000;
    16'b1111111110110001 : data_out = 24'b000000000001110110011111;
    16'b1111111110110010 : data_out = 24'b000000000001110110100111;
    16'b1111111110110011 : data_out = 24'b000000000001110110101110;
    16'b1111111110110100 : data_out = 24'b000000000001110110110110;
    16'b1111111110110101 : data_out = 24'b000000000001110110111101;
    16'b1111111110110110 : data_out = 24'b000000000001110111000100;
    16'b1111111110110111 : data_out = 24'b000000000001110111001100;
    16'b1111111110111000 : data_out = 24'b000000000001110111010011;
    16'b1111111110111001 : data_out = 24'b000000000001110111011011;
    16'b1111111110111010 : data_out = 24'b000000000001110111100010;
    16'b1111111110111011 : data_out = 24'b000000000001110111101010;
    16'b1111111110111100 : data_out = 24'b000000000001110111110001;
    16'b1111111110111101 : data_out = 24'b000000000001110111111001;
    16'b1111111110111110 : data_out = 24'b000000000001111000000000;
    16'b1111111110111111 : data_out = 24'b000000000001111000001000;
    16'b1111111111000000 : data_out = 24'b000000000001111000001111;
    16'b1111111111000001 : data_out = 24'b000000000001111000010111;
    16'b1111111111000010 : data_out = 24'b000000000001111000011110;
    16'b1111111111000011 : data_out = 24'b000000000001111000100110;
    16'b1111111111000100 : data_out = 24'b000000000001111000101101;
    16'b1111111111000101 : data_out = 24'b000000000001111000110101;
    16'b1111111111000110 : data_out = 24'b000000000001111000111100;
    16'b1111111111000111 : data_out = 24'b000000000001111001000100;
    16'b1111111111001000 : data_out = 24'b000000000001111001001100;
    16'b1111111111001001 : data_out = 24'b000000000001111001010011;
    16'b1111111111001010 : data_out = 24'b000000000001111001011011;
    16'b1111111111001011 : data_out = 24'b000000000001111001100010;
    16'b1111111111001100 : data_out = 24'b000000000001111001101010;
    16'b1111111111001101 : data_out = 24'b000000000001111001110001;
    16'b1111111111001110 : data_out = 24'b000000000001111001111001;
    16'b1111111111001111 : data_out = 24'b000000000001111010000001;
    16'b1111111111010000 : data_out = 24'b000000000001111010001000;
    16'b1111111111010001 : data_out = 24'b000000000001111010010000;
    16'b1111111111010010 : data_out = 24'b000000000001111010011000;
    16'b1111111111010011 : data_out = 24'b000000000001111010011111;
    16'b1111111111010100 : data_out = 24'b000000000001111010100111;
    16'b1111111111010101 : data_out = 24'b000000000001111010101111;
    16'b1111111111010110 : data_out = 24'b000000000001111010110110;
    16'b1111111111010111 : data_out = 24'b000000000001111010111110;
    16'b1111111111011000 : data_out = 24'b000000000001111011000110;
    16'b1111111111011001 : data_out = 24'b000000000001111011001101;
    16'b1111111111011010 : data_out = 24'b000000000001111011010101;
    16'b1111111111011011 : data_out = 24'b000000000001111011011101;
    16'b1111111111011100 : data_out = 24'b000000000001111011100101;
    16'b1111111111011101 : data_out = 24'b000000000001111011101100;
    16'b1111111111011110 : data_out = 24'b000000000001111011110100;
    16'b1111111111011111 : data_out = 24'b000000000001111011111100;
    16'b1111111111100000 : data_out = 24'b000000000001111100000011;
    16'b1111111111100001 : data_out = 24'b000000000001111100001011;
    16'b1111111111100010 : data_out = 24'b000000000001111100010011;
    16'b1111111111100011 : data_out = 24'b000000000001111100011011;
    16'b1111111111100100 : data_out = 24'b000000000001111100100011;
    16'b1111111111100101 : data_out = 24'b000000000001111100101010;
    16'b1111111111100110 : data_out = 24'b000000000001111100110010;
    16'b1111111111100111 : data_out = 24'b000000000001111100111010;
    16'b1111111111101000 : data_out = 24'b000000000001111101000010;
    16'b1111111111101001 : data_out = 24'b000000000001111101001010;
    16'b1111111111101010 : data_out = 24'b000000000001111101010001;
    16'b1111111111101011 : data_out = 24'b000000000001111101011001;
    16'b1111111111101100 : data_out = 24'b000000000001111101100001;
    16'b1111111111101101 : data_out = 24'b000000000001111101101001;
    16'b1111111111101110 : data_out = 24'b000000000001111101110001;
    16'b1111111111101111 : data_out = 24'b000000000001111101111001;
    16'b1111111111110000 : data_out = 24'b000000000001111110000000;
    16'b1111111111110001 : data_out = 24'b000000000001111110001000;
    16'b1111111111110010 : data_out = 24'b000000000001111110010000;
    16'b1111111111110011 : data_out = 24'b000000000001111110011000;
    16'b1111111111110100 : data_out = 24'b000000000001111110100000;
    16'b1111111111110101 : data_out = 24'b000000000001111110101000;
    16'b1111111111110110 : data_out = 24'b000000000001111110110000;
    16'b1111111111110111 : data_out = 24'b000000000001111110111000;
    16'b1111111111111000 : data_out = 24'b000000000001111111000000;
    16'b1111111111111001 : data_out = 24'b000000000001111111001000;
    16'b1111111111111010 : data_out = 24'b000000000001111111010000;
    16'b1111111111111011 : data_out = 24'b000000000001111111011000;
    16'b1111111111111100 : data_out = 24'b000000000001111111100000;
    16'b1111111111111101 : data_out = 24'b000000000001111111101000;
    16'b1111111111111110 : data_out = 24'b000000000001111111110000;
    16'b1111111111111111 : data_out = 24'b000000000001111111111000;
    16'b0000000000000000 : data_out = 24'b000000000010000000000000;
    16'b0000000000000001 : data_out = 24'b000000000010000000001000;
    16'b0000000000000010 : data_out = 24'b000000000010000000010000;
    16'b0000000000000011 : data_out = 24'b000000000010000000011000;
    16'b0000000000000100 : data_out = 24'b000000000010000000100000;
    16'b0000000000000101 : data_out = 24'b000000000010000000101000;
    16'b0000000000000110 : data_out = 24'b000000000010000000110000;
    16'b0000000000000111 : data_out = 24'b000000000010000000111000;
    16'b0000000000001000 : data_out = 24'b000000000010000001000000;
    16'b0000000000001001 : data_out = 24'b000000000010000001001000;
    16'b0000000000001010 : data_out = 24'b000000000010000001010000;
    16'b0000000000001011 : data_out = 24'b000000000010000001011000;
    16'b0000000000001100 : data_out = 24'b000000000010000001100000;
    16'b0000000000001101 : data_out = 24'b000000000010000001101000;
    16'b0000000000001110 : data_out = 24'b000000000010000001110000;
    16'b0000000000001111 : data_out = 24'b000000000010000001111000;
    16'b0000000000010000 : data_out = 24'b000000000010000010000001;
    16'b0000000000010001 : data_out = 24'b000000000010000010001001;
    16'b0000000000010010 : data_out = 24'b000000000010000010010001;
    16'b0000000000010011 : data_out = 24'b000000000010000010011001;
    16'b0000000000010100 : data_out = 24'b000000000010000010100001;
    16'b0000000000010101 : data_out = 24'b000000000010000010101001;
    16'b0000000000010110 : data_out = 24'b000000000010000010110001;
    16'b0000000000010111 : data_out = 24'b000000000010000010111010;
    16'b0000000000011000 : data_out = 24'b000000000010000011000010;
    16'b0000000000011001 : data_out = 24'b000000000010000011001010;
    16'b0000000000011010 : data_out = 24'b000000000010000011010010;
    16'b0000000000011011 : data_out = 24'b000000000010000011011010;
    16'b0000000000011100 : data_out = 24'b000000000010000011100011;
    16'b0000000000011101 : data_out = 24'b000000000010000011101011;
    16'b0000000000011110 : data_out = 24'b000000000010000011110011;
    16'b0000000000011111 : data_out = 24'b000000000010000011111011;
    16'b0000000000100000 : data_out = 24'b000000000010000100000100;
    16'b0000000000100001 : data_out = 24'b000000000010000100001100;
    16'b0000000000100010 : data_out = 24'b000000000010000100010100;
    16'b0000000000100011 : data_out = 24'b000000000010000100011100;
    16'b0000000000100100 : data_out = 24'b000000000010000100100101;
    16'b0000000000100101 : data_out = 24'b000000000010000100101101;
    16'b0000000000100110 : data_out = 24'b000000000010000100110101;
    16'b0000000000100111 : data_out = 24'b000000000010000100111110;
    16'b0000000000101000 : data_out = 24'b000000000010000101000110;
    16'b0000000000101001 : data_out = 24'b000000000010000101001110;
    16'b0000000000101010 : data_out = 24'b000000000010000101010110;
    16'b0000000000101011 : data_out = 24'b000000000010000101011111;
    16'b0000000000101100 : data_out = 24'b000000000010000101100111;
    16'b0000000000101101 : data_out = 24'b000000000010000101110000;
    16'b0000000000101110 : data_out = 24'b000000000010000101111000;
    16'b0000000000101111 : data_out = 24'b000000000010000110000000;
    16'b0000000000110000 : data_out = 24'b000000000010000110001001;
    16'b0000000000110001 : data_out = 24'b000000000010000110010001;
    16'b0000000000110010 : data_out = 24'b000000000010000110011001;
    16'b0000000000110011 : data_out = 24'b000000000010000110100010;
    16'b0000000000110100 : data_out = 24'b000000000010000110101010;
    16'b0000000000110101 : data_out = 24'b000000000010000110110011;
    16'b0000000000110110 : data_out = 24'b000000000010000110111011;
    16'b0000000000110111 : data_out = 24'b000000000010000111000100;
    16'b0000000000111000 : data_out = 24'b000000000010000111001100;
    16'b0000000000111001 : data_out = 24'b000000000010000111010100;
    16'b0000000000111010 : data_out = 24'b000000000010000111011101;
    16'b0000000000111011 : data_out = 24'b000000000010000111100101;
    16'b0000000000111100 : data_out = 24'b000000000010000111101110;
    16'b0000000000111101 : data_out = 24'b000000000010000111110110;
    16'b0000000000111110 : data_out = 24'b000000000010000111111111;
    16'b0000000000111111 : data_out = 24'b000000000010001000000111;
    16'b0000000001000000 : data_out = 24'b000000000010001000010000;
    16'b0000000001000001 : data_out = 24'b000000000010001000011000;
    16'b0000000001000010 : data_out = 24'b000000000010001000100001;
    16'b0000000001000011 : data_out = 24'b000000000010001000101001;
    16'b0000000001000100 : data_out = 24'b000000000010001000110010;
    16'b0000000001000101 : data_out = 24'b000000000010001000111011;
    16'b0000000001000110 : data_out = 24'b000000000010001001000011;
    16'b0000000001000111 : data_out = 24'b000000000010001001001100;
    16'b0000000001001000 : data_out = 24'b000000000010001001010100;
    16'b0000000001001001 : data_out = 24'b000000000010001001011101;
    16'b0000000001001010 : data_out = 24'b000000000010001001100101;
    16'b0000000001001011 : data_out = 24'b000000000010001001101110;
    16'b0000000001001100 : data_out = 24'b000000000010001001110111;
    16'b0000000001001101 : data_out = 24'b000000000010001001111111;
    16'b0000000001001110 : data_out = 24'b000000000010001010001000;
    16'b0000000001001111 : data_out = 24'b000000000010001010010001;
    16'b0000000001010000 : data_out = 24'b000000000010001010011001;
    16'b0000000001010001 : data_out = 24'b000000000010001010100010;
    16'b0000000001010010 : data_out = 24'b000000000010001010101010;
    16'b0000000001010011 : data_out = 24'b000000000010001010110011;
    16'b0000000001010100 : data_out = 24'b000000000010001010111100;
    16'b0000000001010101 : data_out = 24'b000000000010001011000101;
    16'b0000000001010110 : data_out = 24'b000000000010001011001101;
    16'b0000000001010111 : data_out = 24'b000000000010001011010110;
    16'b0000000001011000 : data_out = 24'b000000000010001011011111;
    16'b0000000001011001 : data_out = 24'b000000000010001011100111;
    16'b0000000001011010 : data_out = 24'b000000000010001011110000;
    16'b0000000001011011 : data_out = 24'b000000000010001011111001;
    16'b0000000001011100 : data_out = 24'b000000000010001100000010;
    16'b0000000001011101 : data_out = 24'b000000000010001100001010;
    16'b0000000001011110 : data_out = 24'b000000000010001100010011;
    16'b0000000001011111 : data_out = 24'b000000000010001100011100;
    16'b0000000001100000 : data_out = 24'b000000000010001100100101;
    16'b0000000001100001 : data_out = 24'b000000000010001100101101;
    16'b0000000001100010 : data_out = 24'b000000000010001100110110;
    16'b0000000001100011 : data_out = 24'b000000000010001100111111;
    16'b0000000001100100 : data_out = 24'b000000000010001101001000;
    16'b0000000001100101 : data_out = 24'b000000000010001101010001;
    16'b0000000001100110 : data_out = 24'b000000000010001101011010;
    16'b0000000001100111 : data_out = 24'b000000000010001101100010;
    16'b0000000001101000 : data_out = 24'b000000000010001101101011;
    16'b0000000001101001 : data_out = 24'b000000000010001101110100;
    16'b0000000001101010 : data_out = 24'b000000000010001101111101;
    16'b0000000001101011 : data_out = 24'b000000000010001110000110;
    16'b0000000001101100 : data_out = 24'b000000000010001110001111;
    16'b0000000001101101 : data_out = 24'b000000000010001110011000;
    16'b0000000001101110 : data_out = 24'b000000000010001110100001;
    16'b0000000001101111 : data_out = 24'b000000000010001110101001;
    16'b0000000001110000 : data_out = 24'b000000000010001110110010;
    16'b0000000001110001 : data_out = 24'b000000000010001110111011;
    16'b0000000001110010 : data_out = 24'b000000000010001111000100;
    16'b0000000001110011 : data_out = 24'b000000000010001111001101;
    16'b0000000001110100 : data_out = 24'b000000000010001111010110;
    16'b0000000001110101 : data_out = 24'b000000000010001111011111;
    16'b0000000001110110 : data_out = 24'b000000000010001111101000;
    16'b0000000001110111 : data_out = 24'b000000000010001111110001;
    16'b0000000001111000 : data_out = 24'b000000000010001111111010;
    16'b0000000001111001 : data_out = 24'b000000000010010000000011;
    16'b0000000001111010 : data_out = 24'b000000000010010000001100;
    16'b0000000001111011 : data_out = 24'b000000000010010000010101;
    16'b0000000001111100 : data_out = 24'b000000000010010000011110;
    16'b0000000001111101 : data_out = 24'b000000000010010000100111;
    16'b0000000001111110 : data_out = 24'b000000000010010000110000;
    16'b0000000001111111 : data_out = 24'b000000000010010000111001;
    16'b0000000010000000 : data_out = 24'b000000000010010001000010;
    16'b0000000010000001 : data_out = 24'b000000000010010001001011;
    16'b0000000010000010 : data_out = 24'b000000000010010001010100;
    16'b0000000010000011 : data_out = 24'b000000000010010001011101;
    16'b0000000010000100 : data_out = 24'b000000000010010001100111;
    16'b0000000010000101 : data_out = 24'b000000000010010001110000;
    16'b0000000010000110 : data_out = 24'b000000000010010001111001;
    16'b0000000010000111 : data_out = 24'b000000000010010010000010;
    16'b0000000010001000 : data_out = 24'b000000000010010010001011;
    16'b0000000010001001 : data_out = 24'b000000000010010010010100;
    16'b0000000010001010 : data_out = 24'b000000000010010010011101;
    16'b0000000010001011 : data_out = 24'b000000000010010010100111;
    16'b0000000010001100 : data_out = 24'b000000000010010010110000;
    16'b0000000010001101 : data_out = 24'b000000000010010010111001;
    16'b0000000010001110 : data_out = 24'b000000000010010011000010;
    16'b0000000010001111 : data_out = 24'b000000000010010011001011;
    16'b0000000010010000 : data_out = 24'b000000000010010011010100;
    16'b0000000010010001 : data_out = 24'b000000000010010011011110;
    16'b0000000010010010 : data_out = 24'b000000000010010011100111;
    16'b0000000010010011 : data_out = 24'b000000000010010011110000;
    16'b0000000010010100 : data_out = 24'b000000000010010011111001;
    16'b0000000010010101 : data_out = 24'b000000000010010100000011;
    16'b0000000010010110 : data_out = 24'b000000000010010100001100;
    16'b0000000010010111 : data_out = 24'b000000000010010100010101;
    16'b0000000010011000 : data_out = 24'b000000000010010100011110;
    16'b0000000010011001 : data_out = 24'b000000000010010100101000;
    16'b0000000010011010 : data_out = 24'b000000000010010100110001;
    16'b0000000010011011 : data_out = 24'b000000000010010100111010;
    16'b0000000010011100 : data_out = 24'b000000000010010101000100;
    16'b0000000010011101 : data_out = 24'b000000000010010101001101;
    16'b0000000010011110 : data_out = 24'b000000000010010101010110;
    16'b0000000010011111 : data_out = 24'b000000000010010101100000;
    16'b0000000010100000 : data_out = 24'b000000000010010101101001;
    16'b0000000010100001 : data_out = 24'b000000000010010101110010;
    16'b0000000010100010 : data_out = 24'b000000000010010101111100;
    16'b0000000010100011 : data_out = 24'b000000000010010110000101;
    16'b0000000010100100 : data_out = 24'b000000000010010110001110;
    16'b0000000010100101 : data_out = 24'b000000000010010110011000;
    16'b0000000010100110 : data_out = 24'b000000000010010110100001;
    16'b0000000010100111 : data_out = 24'b000000000010010110101011;
    16'b0000000010101000 : data_out = 24'b000000000010010110110100;
    16'b0000000010101001 : data_out = 24'b000000000010010110111101;
    16'b0000000010101010 : data_out = 24'b000000000010010111000111;
    16'b0000000010101011 : data_out = 24'b000000000010010111010000;
    16'b0000000010101100 : data_out = 24'b000000000010010111011010;
    16'b0000000010101101 : data_out = 24'b000000000010010111100011;
    16'b0000000010101110 : data_out = 24'b000000000010010111101101;
    16'b0000000010101111 : data_out = 24'b000000000010010111110110;
    16'b0000000010110000 : data_out = 24'b000000000010011000000000;
    16'b0000000010110001 : data_out = 24'b000000000010011000001001;
    16'b0000000010110010 : data_out = 24'b000000000010011000010011;
    16'b0000000010110011 : data_out = 24'b000000000010011000011100;
    16'b0000000010110100 : data_out = 24'b000000000010011000100110;
    16'b0000000010110101 : data_out = 24'b000000000010011000101111;
    16'b0000000010110110 : data_out = 24'b000000000010011000111001;
    16'b0000000010110111 : data_out = 24'b000000000010011001000010;
    16'b0000000010111000 : data_out = 24'b000000000010011001001100;
    16'b0000000010111001 : data_out = 24'b000000000010011001010110;
    16'b0000000010111010 : data_out = 24'b000000000010011001011111;
    16'b0000000010111011 : data_out = 24'b000000000010011001101001;
    16'b0000000010111100 : data_out = 24'b000000000010011001110010;
    16'b0000000010111101 : data_out = 24'b000000000010011001111100;
    16'b0000000010111110 : data_out = 24'b000000000010011010000110;
    16'b0000000010111111 : data_out = 24'b000000000010011010001111;
    16'b0000000011000000 : data_out = 24'b000000000010011010011001;
    16'b0000000011000001 : data_out = 24'b000000000010011010100011;
    16'b0000000011000010 : data_out = 24'b000000000010011010101100;
    16'b0000000011000011 : data_out = 24'b000000000010011010110110;
    16'b0000000011000100 : data_out = 24'b000000000010011011000000;
    16'b0000000011000101 : data_out = 24'b000000000010011011001001;
    16'b0000000011000110 : data_out = 24'b000000000010011011010011;
    16'b0000000011000111 : data_out = 24'b000000000010011011011101;
    16'b0000000011001000 : data_out = 24'b000000000010011011100110;
    16'b0000000011001001 : data_out = 24'b000000000010011011110000;
    16'b0000000011001010 : data_out = 24'b000000000010011011111010;
    16'b0000000011001011 : data_out = 24'b000000000010011100000100;
    16'b0000000011001100 : data_out = 24'b000000000010011100001101;
    16'b0000000011001101 : data_out = 24'b000000000010011100010111;
    16'b0000000011001110 : data_out = 24'b000000000010011100100001;
    16'b0000000011001111 : data_out = 24'b000000000010011100101011;
    16'b0000000011010000 : data_out = 24'b000000000010011100110101;
    16'b0000000011010001 : data_out = 24'b000000000010011100111110;
    16'b0000000011010010 : data_out = 24'b000000000010011101001000;
    16'b0000000011010011 : data_out = 24'b000000000010011101010010;
    16'b0000000011010100 : data_out = 24'b000000000010011101011100;
    16'b0000000011010101 : data_out = 24'b000000000010011101100110;
    16'b0000000011010110 : data_out = 24'b000000000010011101110000;
    16'b0000000011010111 : data_out = 24'b000000000010011101111001;
    16'b0000000011011000 : data_out = 24'b000000000010011110000011;
    16'b0000000011011001 : data_out = 24'b000000000010011110001101;
    16'b0000000011011010 : data_out = 24'b000000000010011110010111;
    16'b0000000011011011 : data_out = 24'b000000000010011110100001;
    16'b0000000011011100 : data_out = 24'b000000000010011110101011;
    16'b0000000011011101 : data_out = 24'b000000000010011110110101;
    16'b0000000011011110 : data_out = 24'b000000000010011110111111;
    16'b0000000011011111 : data_out = 24'b000000000010011111001001;
    16'b0000000011100000 : data_out = 24'b000000000010011111010011;
    16'b0000000011100001 : data_out = 24'b000000000010011111011101;
    16'b0000000011100010 : data_out = 24'b000000000010011111100111;
    16'b0000000011100011 : data_out = 24'b000000000010011111110001;
    16'b0000000011100100 : data_out = 24'b000000000010011111111011;
    16'b0000000011100101 : data_out = 24'b000000000010100000000101;
    16'b0000000011100110 : data_out = 24'b000000000010100000001111;
    16'b0000000011100111 : data_out = 24'b000000000010100000011001;
    16'b0000000011101000 : data_out = 24'b000000000010100000100011;
    16'b0000000011101001 : data_out = 24'b000000000010100000101101;
    16'b0000000011101010 : data_out = 24'b000000000010100000110111;
    16'b0000000011101011 : data_out = 24'b000000000010100001000001;
    16'b0000000011101100 : data_out = 24'b000000000010100001001011;
    16'b0000000011101101 : data_out = 24'b000000000010100001010101;
    16'b0000000011101110 : data_out = 24'b000000000010100001011111;
    16'b0000000011101111 : data_out = 24'b000000000010100001101001;
    16'b0000000011110000 : data_out = 24'b000000000010100001110011;
    16'b0000000011110001 : data_out = 24'b000000000010100001111101;
    16'b0000000011110010 : data_out = 24'b000000000010100010000111;
    16'b0000000011110011 : data_out = 24'b000000000010100010010010;
    16'b0000000011110100 : data_out = 24'b000000000010100010011100;
    16'b0000000011110101 : data_out = 24'b000000000010100010100110;
    16'b0000000011110110 : data_out = 24'b000000000010100010110000;
    16'b0000000011110111 : data_out = 24'b000000000010100010111010;
    16'b0000000011111000 : data_out = 24'b000000000010100011000100;
    16'b0000000011111001 : data_out = 24'b000000000010100011001111;
    16'b0000000011111010 : data_out = 24'b000000000010100011011001;
    16'b0000000011111011 : data_out = 24'b000000000010100011100011;
    16'b0000000011111100 : data_out = 24'b000000000010100011101101;
    16'b0000000011111101 : data_out = 24'b000000000010100011110111;
    16'b0000000011111110 : data_out = 24'b000000000010100100000010;
    16'b0000000011111111 : data_out = 24'b000000000010100100001100;
    16'b0000000100000000 : data_out = 24'b000000000010100100010110;
    16'b0000000100000001 : data_out = 24'b000000000010100100100001;
    16'b0000000100000010 : data_out = 24'b000000000010100100101011;
    16'b0000000100000011 : data_out = 24'b000000000010100100110101;
    16'b0000000100000100 : data_out = 24'b000000000010100100111111;
    16'b0000000100000101 : data_out = 24'b000000000010100101001010;
    16'b0000000100000110 : data_out = 24'b000000000010100101010100;
    16'b0000000100000111 : data_out = 24'b000000000010100101011110;
    16'b0000000100001000 : data_out = 24'b000000000010100101101001;
    16'b0000000100001001 : data_out = 24'b000000000010100101110011;
    16'b0000000100001010 : data_out = 24'b000000000010100101111101;
    16'b0000000100001011 : data_out = 24'b000000000010100110001000;
    16'b0000000100001100 : data_out = 24'b000000000010100110010010;
    16'b0000000100001101 : data_out = 24'b000000000010100110011101;
    16'b0000000100001110 : data_out = 24'b000000000010100110100111;
    16'b0000000100001111 : data_out = 24'b000000000010100110110001;
    16'b0000000100010000 : data_out = 24'b000000000010100110111100;
    16'b0000000100010001 : data_out = 24'b000000000010100111000110;
    16'b0000000100010010 : data_out = 24'b000000000010100111010001;
    16'b0000000100010011 : data_out = 24'b000000000010100111011011;
    16'b0000000100010100 : data_out = 24'b000000000010100111100110;
    16'b0000000100010101 : data_out = 24'b000000000010100111110000;
    16'b0000000100010110 : data_out = 24'b000000000010100111111011;
    16'b0000000100010111 : data_out = 24'b000000000010101000000101;
    16'b0000000100011000 : data_out = 24'b000000000010101000010000;
    16'b0000000100011001 : data_out = 24'b000000000010101000011010;
    16'b0000000100011010 : data_out = 24'b000000000010101000100101;
    16'b0000000100011011 : data_out = 24'b000000000010101000101111;
    16'b0000000100011100 : data_out = 24'b000000000010101000111010;
    16'b0000000100011101 : data_out = 24'b000000000010101001000100;
    16'b0000000100011110 : data_out = 24'b000000000010101001001111;
    16'b0000000100011111 : data_out = 24'b000000000010101001011010;
    16'b0000000100100000 : data_out = 24'b000000000010101001100100;
    16'b0000000100100001 : data_out = 24'b000000000010101001101111;
    16'b0000000100100010 : data_out = 24'b000000000010101001111001;
    16'b0000000100100011 : data_out = 24'b000000000010101010000100;
    16'b0000000100100100 : data_out = 24'b000000000010101010001111;
    16'b0000000100100101 : data_out = 24'b000000000010101010011001;
    16'b0000000100100110 : data_out = 24'b000000000010101010100100;
    16'b0000000100100111 : data_out = 24'b000000000010101010101111;
    16'b0000000100101000 : data_out = 24'b000000000010101010111001;
    16'b0000000100101001 : data_out = 24'b000000000010101011000100;
    16'b0000000100101010 : data_out = 24'b000000000010101011001111;
    16'b0000000100101011 : data_out = 24'b000000000010101011011001;
    16'b0000000100101100 : data_out = 24'b000000000010101011100100;
    16'b0000000100101101 : data_out = 24'b000000000010101011101111;
    16'b0000000100101110 : data_out = 24'b000000000010101011111010;
    16'b0000000100101111 : data_out = 24'b000000000010101100000100;
    16'b0000000100110000 : data_out = 24'b000000000010101100001111;
    16'b0000000100110001 : data_out = 24'b000000000010101100011010;
    16'b0000000100110010 : data_out = 24'b000000000010101100100101;
    16'b0000000100110011 : data_out = 24'b000000000010101100101111;
    16'b0000000100110100 : data_out = 24'b000000000010101100111010;
    16'b0000000100110101 : data_out = 24'b000000000010101101000101;
    16'b0000000100110110 : data_out = 24'b000000000010101101010000;
    16'b0000000100110111 : data_out = 24'b000000000010101101011011;
    16'b0000000100111000 : data_out = 24'b000000000010101101100101;
    16'b0000000100111001 : data_out = 24'b000000000010101101110000;
    16'b0000000100111010 : data_out = 24'b000000000010101101111011;
    16'b0000000100111011 : data_out = 24'b000000000010101110000110;
    16'b0000000100111100 : data_out = 24'b000000000010101110010001;
    16'b0000000100111101 : data_out = 24'b000000000010101110011100;
    16'b0000000100111110 : data_out = 24'b000000000010101110100111;
    16'b0000000100111111 : data_out = 24'b000000000010101110110010;
    16'b0000000101000000 : data_out = 24'b000000000010101110111101;
    16'b0000000101000001 : data_out = 24'b000000000010101111001000;
    16'b0000000101000010 : data_out = 24'b000000000010101111010011;
    16'b0000000101000011 : data_out = 24'b000000000010101111011101;
    16'b0000000101000100 : data_out = 24'b000000000010101111101000;
    16'b0000000101000101 : data_out = 24'b000000000010101111110011;
    16'b0000000101000110 : data_out = 24'b000000000010101111111110;
    16'b0000000101000111 : data_out = 24'b000000000010110000001001;
    16'b0000000101001000 : data_out = 24'b000000000010110000010100;
    16'b0000000101001001 : data_out = 24'b000000000010110000011111;
    16'b0000000101001010 : data_out = 24'b000000000010110000101011;
    16'b0000000101001011 : data_out = 24'b000000000010110000110110;
    16'b0000000101001100 : data_out = 24'b000000000010110001000001;
    16'b0000000101001101 : data_out = 24'b000000000010110001001100;
    16'b0000000101001110 : data_out = 24'b000000000010110001010111;
    16'b0000000101001111 : data_out = 24'b000000000010110001100010;
    16'b0000000101010000 : data_out = 24'b000000000010110001101101;
    16'b0000000101010001 : data_out = 24'b000000000010110001111000;
    16'b0000000101010010 : data_out = 24'b000000000010110010000011;
    16'b0000000101010011 : data_out = 24'b000000000010110010001110;
    16'b0000000101010100 : data_out = 24'b000000000010110010011001;
    16'b0000000101010101 : data_out = 24'b000000000010110010100101;
    16'b0000000101010110 : data_out = 24'b000000000010110010110000;
    16'b0000000101010111 : data_out = 24'b000000000010110010111011;
    16'b0000000101011000 : data_out = 24'b000000000010110011000110;
    16'b0000000101011001 : data_out = 24'b000000000010110011010001;
    16'b0000000101011010 : data_out = 24'b000000000010110011011101;
    16'b0000000101011011 : data_out = 24'b000000000010110011101000;
    16'b0000000101011100 : data_out = 24'b000000000010110011110011;
    16'b0000000101011101 : data_out = 24'b000000000010110011111110;
    16'b0000000101011110 : data_out = 24'b000000000010110100001010;
    16'b0000000101011111 : data_out = 24'b000000000010110100010101;
    16'b0000000101100000 : data_out = 24'b000000000010110100100000;
    16'b0000000101100001 : data_out = 24'b000000000010110100101011;
    16'b0000000101100010 : data_out = 24'b000000000010110100110111;
    16'b0000000101100011 : data_out = 24'b000000000010110101000010;
    16'b0000000101100100 : data_out = 24'b000000000010110101001101;
    16'b0000000101100101 : data_out = 24'b000000000010110101011001;
    16'b0000000101100110 : data_out = 24'b000000000010110101100100;
    16'b0000000101100111 : data_out = 24'b000000000010110101101111;
    16'b0000000101101000 : data_out = 24'b000000000010110101111011;
    16'b0000000101101001 : data_out = 24'b000000000010110110000110;
    16'b0000000101101010 : data_out = 24'b000000000010110110010001;
    16'b0000000101101011 : data_out = 24'b000000000010110110011101;
    16'b0000000101101100 : data_out = 24'b000000000010110110101000;
    16'b0000000101101101 : data_out = 24'b000000000010110110110100;
    16'b0000000101101110 : data_out = 24'b000000000010110110111111;
    16'b0000000101101111 : data_out = 24'b000000000010110111001011;
    16'b0000000101110000 : data_out = 24'b000000000010110111010110;
    16'b0000000101110001 : data_out = 24'b000000000010110111100001;
    16'b0000000101110010 : data_out = 24'b000000000010110111101101;
    16'b0000000101110011 : data_out = 24'b000000000010110111111000;
    16'b0000000101110100 : data_out = 24'b000000000010111000000100;
    16'b0000000101110101 : data_out = 24'b000000000010111000001111;
    16'b0000000101110110 : data_out = 24'b000000000010111000011011;
    16'b0000000101110111 : data_out = 24'b000000000010111000100110;
    16'b0000000101111000 : data_out = 24'b000000000010111000110010;
    16'b0000000101111001 : data_out = 24'b000000000010111000111110;
    16'b0000000101111010 : data_out = 24'b000000000010111001001001;
    16'b0000000101111011 : data_out = 24'b000000000010111001010101;
    16'b0000000101111100 : data_out = 24'b000000000010111001100000;
    16'b0000000101111101 : data_out = 24'b000000000010111001101100;
    16'b0000000101111110 : data_out = 24'b000000000010111001111000;
    16'b0000000101111111 : data_out = 24'b000000000010111010000011;
    16'b0000000110000000 : data_out = 24'b000000000010111010001111;
    16'b0000000110000001 : data_out = 24'b000000000010111010011010;
    16'b0000000110000010 : data_out = 24'b000000000010111010100110;
    16'b0000000110000011 : data_out = 24'b000000000010111010110010;
    16'b0000000110000100 : data_out = 24'b000000000010111010111101;
    16'b0000000110000101 : data_out = 24'b000000000010111011001001;
    16'b0000000110000110 : data_out = 24'b000000000010111011010101;
    16'b0000000110000111 : data_out = 24'b000000000010111011100001;
    16'b0000000110001000 : data_out = 24'b000000000010111011101100;
    16'b0000000110001001 : data_out = 24'b000000000010111011111000;
    16'b0000000110001010 : data_out = 24'b000000000010111100000100;
    16'b0000000110001011 : data_out = 24'b000000000010111100010000;
    16'b0000000110001100 : data_out = 24'b000000000010111100011011;
    16'b0000000110001101 : data_out = 24'b000000000010111100100111;
    16'b0000000110001110 : data_out = 24'b000000000010111100110011;
    16'b0000000110001111 : data_out = 24'b000000000010111100111111;
    16'b0000000110010000 : data_out = 24'b000000000010111101001010;
    16'b0000000110010001 : data_out = 24'b000000000010111101010110;
    16'b0000000110010010 : data_out = 24'b000000000010111101100010;
    16'b0000000110010011 : data_out = 24'b000000000010111101101110;
    16'b0000000110010100 : data_out = 24'b000000000010111101111010;
    16'b0000000110010101 : data_out = 24'b000000000010111110000110;
    16'b0000000110010110 : data_out = 24'b000000000010111110010010;
    16'b0000000110010111 : data_out = 24'b000000000010111110011110;
    16'b0000000110011000 : data_out = 24'b000000000010111110101001;
    16'b0000000110011001 : data_out = 24'b000000000010111110110101;
    16'b0000000110011010 : data_out = 24'b000000000010111111000001;
    16'b0000000110011011 : data_out = 24'b000000000010111111001101;
    16'b0000000110011100 : data_out = 24'b000000000010111111011001;
    16'b0000000110011101 : data_out = 24'b000000000010111111100101;
    16'b0000000110011110 : data_out = 24'b000000000010111111110001;
    16'b0000000110011111 : data_out = 24'b000000000010111111111101;
    16'b0000000110100000 : data_out = 24'b000000000011000000001001;
    16'b0000000110100001 : data_out = 24'b000000000011000000010101;
    16'b0000000110100010 : data_out = 24'b000000000011000000100001;
    16'b0000000110100011 : data_out = 24'b000000000011000000101101;
    16'b0000000110100100 : data_out = 24'b000000000011000000111001;
    16'b0000000110100101 : data_out = 24'b000000000011000001000101;
    16'b0000000110100110 : data_out = 24'b000000000011000001010001;
    16'b0000000110100111 : data_out = 24'b000000000011000001011110;
    16'b0000000110101000 : data_out = 24'b000000000011000001101010;
    16'b0000000110101001 : data_out = 24'b000000000011000001110110;
    16'b0000000110101010 : data_out = 24'b000000000011000010000010;
    16'b0000000110101011 : data_out = 24'b000000000011000010001110;
    16'b0000000110101100 : data_out = 24'b000000000011000010011010;
    16'b0000000110101101 : data_out = 24'b000000000011000010100110;
    16'b0000000110101110 : data_out = 24'b000000000011000010110010;
    16'b0000000110101111 : data_out = 24'b000000000011000010111111;
    16'b0000000110110000 : data_out = 24'b000000000011000011001011;
    16'b0000000110110001 : data_out = 24'b000000000011000011010111;
    16'b0000000110110010 : data_out = 24'b000000000011000011100011;
    16'b0000000110110011 : data_out = 24'b000000000011000011101111;
    16'b0000000110110100 : data_out = 24'b000000000011000011111100;
    16'b0000000110110101 : data_out = 24'b000000000011000100001000;
    16'b0000000110110110 : data_out = 24'b000000000011000100010100;
    16'b0000000110110111 : data_out = 24'b000000000011000100100000;
    16'b0000000110111000 : data_out = 24'b000000000011000100101101;
    16'b0000000110111001 : data_out = 24'b000000000011000100111001;
    16'b0000000110111010 : data_out = 24'b000000000011000101000101;
    16'b0000000110111011 : data_out = 24'b000000000011000101010010;
    16'b0000000110111100 : data_out = 24'b000000000011000101011110;
    16'b0000000110111101 : data_out = 24'b000000000011000101101010;
    16'b0000000110111110 : data_out = 24'b000000000011000101110111;
    16'b0000000110111111 : data_out = 24'b000000000011000110000011;
    16'b0000000111000000 : data_out = 24'b000000000011000110010000;
    16'b0000000111000001 : data_out = 24'b000000000011000110011100;
    16'b0000000111000010 : data_out = 24'b000000000011000110101000;
    16'b0000000111000011 : data_out = 24'b000000000011000110110101;
    16'b0000000111000100 : data_out = 24'b000000000011000111000001;
    16'b0000000111000101 : data_out = 24'b000000000011000111001110;
    16'b0000000111000110 : data_out = 24'b000000000011000111011010;
    16'b0000000111000111 : data_out = 24'b000000000011000111100111;
    16'b0000000111001000 : data_out = 24'b000000000011000111110011;
    16'b0000000111001001 : data_out = 24'b000000000011001000000000;
    16'b0000000111001010 : data_out = 24'b000000000011001000001100;
    16'b0000000111001011 : data_out = 24'b000000000011001000011001;
    16'b0000000111001100 : data_out = 24'b000000000011001000100101;
    16'b0000000111001101 : data_out = 24'b000000000011001000110010;
    16'b0000000111001110 : data_out = 24'b000000000011001000111110;
    16'b0000000111001111 : data_out = 24'b000000000011001001001011;
    16'b0000000111010000 : data_out = 24'b000000000011001001010111;
    16'b0000000111010001 : data_out = 24'b000000000011001001100100;
    16'b0000000111010010 : data_out = 24'b000000000011001001110001;
    16'b0000000111010011 : data_out = 24'b000000000011001001111101;
    16'b0000000111010100 : data_out = 24'b000000000011001010001010;
    16'b0000000111010101 : data_out = 24'b000000000011001010010110;
    16'b0000000111010110 : data_out = 24'b000000000011001010100011;
    16'b0000000111010111 : data_out = 24'b000000000011001010110000;
    16'b0000000111011000 : data_out = 24'b000000000011001010111100;
    16'b0000000111011001 : data_out = 24'b000000000011001011001001;
    16'b0000000111011010 : data_out = 24'b000000000011001011010110;
    16'b0000000111011011 : data_out = 24'b000000000011001011100011;
    16'b0000000111011100 : data_out = 24'b000000000011001011101111;
    16'b0000000111011101 : data_out = 24'b000000000011001011111100;
    16'b0000000111011110 : data_out = 24'b000000000011001100001001;
    16'b0000000111011111 : data_out = 24'b000000000011001100010110;
    16'b0000000111100000 : data_out = 24'b000000000011001100100010;
    16'b0000000111100001 : data_out = 24'b000000000011001100101111;
    16'b0000000111100010 : data_out = 24'b000000000011001100111100;
    16'b0000000111100011 : data_out = 24'b000000000011001101001001;
    16'b0000000111100100 : data_out = 24'b000000000011001101010110;
    16'b0000000111100101 : data_out = 24'b000000000011001101100010;
    16'b0000000111100110 : data_out = 24'b000000000011001101101111;
    16'b0000000111100111 : data_out = 24'b000000000011001101111100;
    16'b0000000111101000 : data_out = 24'b000000000011001110001001;
    16'b0000000111101001 : data_out = 24'b000000000011001110010110;
    16'b0000000111101010 : data_out = 24'b000000000011001110100011;
    16'b0000000111101011 : data_out = 24'b000000000011001110110000;
    16'b0000000111101100 : data_out = 24'b000000000011001110111101;
    16'b0000000111101101 : data_out = 24'b000000000011001111001010;
    16'b0000000111101110 : data_out = 24'b000000000011001111010110;
    16'b0000000111101111 : data_out = 24'b000000000011001111100011;
    16'b0000000111110000 : data_out = 24'b000000000011001111110000;
    16'b0000000111110001 : data_out = 24'b000000000011001111111101;
    16'b0000000111110010 : data_out = 24'b000000000011010000001010;
    16'b0000000111110011 : data_out = 24'b000000000011010000010111;
    16'b0000000111110100 : data_out = 24'b000000000011010000100100;
    16'b0000000111110101 : data_out = 24'b000000000011010000110010;
    16'b0000000111110110 : data_out = 24'b000000000011010000111111;
    16'b0000000111110111 : data_out = 24'b000000000011010001001100;
    16'b0000000111111000 : data_out = 24'b000000000011010001011001;
    16'b0000000111111001 : data_out = 24'b000000000011010001100110;
    16'b0000000111111010 : data_out = 24'b000000000011010001110011;
    16'b0000000111111011 : data_out = 24'b000000000011010010000000;
    16'b0000000111111100 : data_out = 24'b000000000011010010001101;
    16'b0000000111111101 : data_out = 24'b000000000011010010011010;
    16'b0000000111111110 : data_out = 24'b000000000011010010100111;
    16'b0000000111111111 : data_out = 24'b000000000011010010110101;
    16'b0000001000000000 : data_out = 24'b000000000011010011000010;
    16'b0000001000000001 : data_out = 24'b000000000011010011001111;
    16'b0000001000000010 : data_out = 24'b000000000011010011011100;
    16'b0000001000000011 : data_out = 24'b000000000011010011101001;
    16'b0000001000000100 : data_out = 24'b000000000011010011110111;
    16'b0000001000000101 : data_out = 24'b000000000011010100000100;
    16'b0000001000000110 : data_out = 24'b000000000011010100010001;
    16'b0000001000000111 : data_out = 24'b000000000011010100011110;
    16'b0000001000001000 : data_out = 24'b000000000011010100101100;
    16'b0000001000001001 : data_out = 24'b000000000011010100111001;
    16'b0000001000001010 : data_out = 24'b000000000011010101000110;
    16'b0000001000001011 : data_out = 24'b000000000011010101010100;
    16'b0000001000001100 : data_out = 24'b000000000011010101100001;
    16'b0000001000001101 : data_out = 24'b000000000011010101101110;
    16'b0000001000001110 : data_out = 24'b000000000011010101111100;
    16'b0000001000001111 : data_out = 24'b000000000011010110001001;
    16'b0000001000010000 : data_out = 24'b000000000011010110010111;
    16'b0000001000010001 : data_out = 24'b000000000011010110100100;
    16'b0000001000010010 : data_out = 24'b000000000011010110110001;
    16'b0000001000010011 : data_out = 24'b000000000011010110111111;
    16'b0000001000010100 : data_out = 24'b000000000011010111001100;
    16'b0000001000010101 : data_out = 24'b000000000011010111011010;
    16'b0000001000010110 : data_out = 24'b000000000011010111100111;
    16'b0000001000010111 : data_out = 24'b000000000011010111110101;
    16'b0000001000011000 : data_out = 24'b000000000011011000000010;
    16'b0000001000011001 : data_out = 24'b000000000011011000010000;
    16'b0000001000011010 : data_out = 24'b000000000011011000011101;
    16'b0000001000011011 : data_out = 24'b000000000011011000101011;
    16'b0000001000011100 : data_out = 24'b000000000011011000111000;
    16'b0000001000011101 : data_out = 24'b000000000011011001000110;
    16'b0000001000011110 : data_out = 24'b000000000011011001010011;
    16'b0000001000011111 : data_out = 24'b000000000011011001100001;
    16'b0000001000100000 : data_out = 24'b000000000011011001101111;
    16'b0000001000100001 : data_out = 24'b000000000011011001111100;
    16'b0000001000100010 : data_out = 24'b000000000011011010001010;
    16'b0000001000100011 : data_out = 24'b000000000011011010010111;
    16'b0000001000100100 : data_out = 24'b000000000011011010100101;
    16'b0000001000100101 : data_out = 24'b000000000011011010110011;
    16'b0000001000100110 : data_out = 24'b000000000011011011000000;
    16'b0000001000100111 : data_out = 24'b000000000011011011001110;
    16'b0000001000101000 : data_out = 24'b000000000011011011011100;
    16'b0000001000101001 : data_out = 24'b000000000011011011101010;
    16'b0000001000101010 : data_out = 24'b000000000011011011110111;
    16'b0000001000101011 : data_out = 24'b000000000011011100000101;
    16'b0000001000101100 : data_out = 24'b000000000011011100010011;
    16'b0000001000101101 : data_out = 24'b000000000011011100100001;
    16'b0000001000101110 : data_out = 24'b000000000011011100101110;
    16'b0000001000101111 : data_out = 24'b000000000011011100111100;
    16'b0000001000110000 : data_out = 24'b000000000011011101001010;
    16'b0000001000110001 : data_out = 24'b000000000011011101011000;
    16'b0000001000110010 : data_out = 24'b000000000011011101100110;
    16'b0000001000110011 : data_out = 24'b000000000011011101110100;
    16'b0000001000110100 : data_out = 24'b000000000011011110000001;
    16'b0000001000110101 : data_out = 24'b000000000011011110001111;
    16'b0000001000110110 : data_out = 24'b000000000011011110011101;
    16'b0000001000110111 : data_out = 24'b000000000011011110101011;
    16'b0000001000111000 : data_out = 24'b000000000011011110111001;
    16'b0000001000111001 : data_out = 24'b000000000011011111000111;
    16'b0000001000111010 : data_out = 24'b000000000011011111010101;
    16'b0000001000111011 : data_out = 24'b000000000011011111100011;
    16'b0000001000111100 : data_out = 24'b000000000011011111110001;
    16'b0000001000111101 : data_out = 24'b000000000011011111111111;
    16'b0000001000111110 : data_out = 24'b000000000011100000001101;
    16'b0000001000111111 : data_out = 24'b000000000011100000011011;
    16'b0000001001000000 : data_out = 24'b000000000011100000101001;
    16'b0000001001000001 : data_out = 24'b000000000011100000110111;
    16'b0000001001000010 : data_out = 24'b000000000011100001000101;
    16'b0000001001000011 : data_out = 24'b000000000011100001010011;
    16'b0000001001000100 : data_out = 24'b000000000011100001100001;
    16'b0000001001000101 : data_out = 24'b000000000011100001101111;
    16'b0000001001000110 : data_out = 24'b000000000011100001111101;
    16'b0000001001000111 : data_out = 24'b000000000011100010001100;
    16'b0000001001001000 : data_out = 24'b000000000011100010011010;
    16'b0000001001001001 : data_out = 24'b000000000011100010101000;
    16'b0000001001001010 : data_out = 24'b000000000011100010110110;
    16'b0000001001001011 : data_out = 24'b000000000011100011000100;
    16'b0000001001001100 : data_out = 24'b000000000011100011010010;
    16'b0000001001001101 : data_out = 24'b000000000011100011100001;
    16'b0000001001001110 : data_out = 24'b000000000011100011101111;
    16'b0000001001001111 : data_out = 24'b000000000011100011111101;
    16'b0000001001010000 : data_out = 24'b000000000011100100001011;
    16'b0000001001010001 : data_out = 24'b000000000011100100011010;
    16'b0000001001010010 : data_out = 24'b000000000011100100101000;
    16'b0000001001010011 : data_out = 24'b000000000011100100110110;
    16'b0000001001010100 : data_out = 24'b000000000011100101000100;
    16'b0000001001010101 : data_out = 24'b000000000011100101010011;
    16'b0000001001010110 : data_out = 24'b000000000011100101100001;
    16'b0000001001010111 : data_out = 24'b000000000011100101101111;
    16'b0000001001011000 : data_out = 24'b000000000011100101111110;
    16'b0000001001011001 : data_out = 24'b000000000011100110001100;
    16'b0000001001011010 : data_out = 24'b000000000011100110011011;
    16'b0000001001011011 : data_out = 24'b000000000011100110101001;
    16'b0000001001011100 : data_out = 24'b000000000011100110110111;
    16'b0000001001011101 : data_out = 24'b000000000011100111000110;
    16'b0000001001011110 : data_out = 24'b000000000011100111010100;
    16'b0000001001011111 : data_out = 24'b000000000011100111100011;
    16'b0000001001100000 : data_out = 24'b000000000011100111110001;
    16'b0000001001100001 : data_out = 24'b000000000011101000000000;
    16'b0000001001100010 : data_out = 24'b000000000011101000001110;
    16'b0000001001100011 : data_out = 24'b000000000011101000011101;
    16'b0000001001100100 : data_out = 24'b000000000011101000101011;
    16'b0000001001100101 : data_out = 24'b000000000011101000111010;
    16'b0000001001100110 : data_out = 24'b000000000011101001001000;
    16'b0000001001100111 : data_out = 24'b000000000011101001010111;
    16'b0000001001101000 : data_out = 24'b000000000011101001100110;
    16'b0000001001101001 : data_out = 24'b000000000011101001110100;
    16'b0000001001101010 : data_out = 24'b000000000011101010000011;
    16'b0000001001101011 : data_out = 24'b000000000011101010010010;
    16'b0000001001101100 : data_out = 24'b000000000011101010100000;
    16'b0000001001101101 : data_out = 24'b000000000011101010101111;
    16'b0000001001101110 : data_out = 24'b000000000011101010111101;
    16'b0000001001101111 : data_out = 24'b000000000011101011001100;
    16'b0000001001110000 : data_out = 24'b000000000011101011011011;
    16'b0000001001110001 : data_out = 24'b000000000011101011101010;
    16'b0000001001110010 : data_out = 24'b000000000011101011111000;
    16'b0000001001110011 : data_out = 24'b000000000011101100000111;
    16'b0000001001110100 : data_out = 24'b000000000011101100010110;
    16'b0000001001110101 : data_out = 24'b000000000011101100100101;
    16'b0000001001110110 : data_out = 24'b000000000011101100110011;
    16'b0000001001110111 : data_out = 24'b000000000011101101000010;
    16'b0000001001111000 : data_out = 24'b000000000011101101010001;
    16'b0000001001111001 : data_out = 24'b000000000011101101100000;
    16'b0000001001111010 : data_out = 24'b000000000011101101101111;
    16'b0000001001111011 : data_out = 24'b000000000011101101111110;
    16'b0000001001111100 : data_out = 24'b000000000011101110001101;
    16'b0000001001111101 : data_out = 24'b000000000011101110011011;
    16'b0000001001111110 : data_out = 24'b000000000011101110101010;
    16'b0000001001111111 : data_out = 24'b000000000011101110111001;
    16'b0000001010000000 : data_out = 24'b000000000011101111001000;
    16'b0000001010000001 : data_out = 24'b000000000011101111010111;
    16'b0000001010000010 : data_out = 24'b000000000011101111100110;
    16'b0000001010000011 : data_out = 24'b000000000011101111110101;
    16'b0000001010000100 : data_out = 24'b000000000011110000000100;
    16'b0000001010000101 : data_out = 24'b000000000011110000010011;
    16'b0000001010000110 : data_out = 24'b000000000011110000100010;
    16'b0000001010000111 : data_out = 24'b000000000011110000110001;
    16'b0000001010001000 : data_out = 24'b000000000011110001000000;
    16'b0000001010001001 : data_out = 24'b000000000011110001001111;
    16'b0000001010001010 : data_out = 24'b000000000011110001011110;
    16'b0000001010001011 : data_out = 24'b000000000011110001101101;
    16'b0000001010001100 : data_out = 24'b000000000011110001111101;
    16'b0000001010001101 : data_out = 24'b000000000011110010001100;
    16'b0000001010001110 : data_out = 24'b000000000011110010011011;
    16'b0000001010001111 : data_out = 24'b000000000011110010101010;
    16'b0000001010010000 : data_out = 24'b000000000011110010111001;
    16'b0000001010010001 : data_out = 24'b000000000011110011001000;
    16'b0000001010010010 : data_out = 24'b000000000011110011011000;
    16'b0000001010010011 : data_out = 24'b000000000011110011100111;
    16'b0000001010010100 : data_out = 24'b000000000011110011110110;
    16'b0000001010010101 : data_out = 24'b000000000011110100000101;
    16'b0000001010010110 : data_out = 24'b000000000011110100010101;
    16'b0000001010010111 : data_out = 24'b000000000011110100100100;
    16'b0000001010011000 : data_out = 24'b000000000011110100110011;
    16'b0000001010011001 : data_out = 24'b000000000011110101000010;
    16'b0000001010011010 : data_out = 24'b000000000011110101010010;
    16'b0000001010011011 : data_out = 24'b000000000011110101100001;
    16'b0000001010011100 : data_out = 24'b000000000011110101110000;
    16'b0000001010011101 : data_out = 24'b000000000011110110000000;
    16'b0000001010011110 : data_out = 24'b000000000011110110001111;
    16'b0000001010011111 : data_out = 24'b000000000011110110011111;
    16'b0000001010100000 : data_out = 24'b000000000011110110101110;
    16'b0000001010100001 : data_out = 24'b000000000011110110111101;
    16'b0000001010100010 : data_out = 24'b000000000011110111001101;
    16'b0000001010100011 : data_out = 24'b000000000011110111011100;
    16'b0000001010100100 : data_out = 24'b000000000011110111101100;
    16'b0000001010100101 : data_out = 24'b000000000011110111111011;
    16'b0000001010100110 : data_out = 24'b000000000011111000001011;
    16'b0000001010100111 : data_out = 24'b000000000011111000011010;
    16'b0000001010101000 : data_out = 24'b000000000011111000101010;
    16'b0000001010101001 : data_out = 24'b000000000011111000111001;
    16'b0000001010101010 : data_out = 24'b000000000011111001001001;
    16'b0000001010101011 : data_out = 24'b000000000011111001011001;
    16'b0000001010101100 : data_out = 24'b000000000011111001101000;
    16'b0000001010101101 : data_out = 24'b000000000011111001111000;
    16'b0000001010101110 : data_out = 24'b000000000011111010000111;
    16'b0000001010101111 : data_out = 24'b000000000011111010010111;
    16'b0000001010110000 : data_out = 24'b000000000011111010100111;
    16'b0000001010110001 : data_out = 24'b000000000011111010110110;
    16'b0000001010110010 : data_out = 24'b000000000011111011000110;
    16'b0000001010110011 : data_out = 24'b000000000011111011010110;
    16'b0000001010110100 : data_out = 24'b000000000011111011100101;
    16'b0000001010110101 : data_out = 24'b000000000011111011110101;
    16'b0000001010110110 : data_out = 24'b000000000011111100000101;
    16'b0000001010110111 : data_out = 24'b000000000011111100010101;
    16'b0000001010111000 : data_out = 24'b000000000011111100100100;
    16'b0000001010111001 : data_out = 24'b000000000011111100110100;
    16'b0000001010111010 : data_out = 24'b000000000011111101000100;
    16'b0000001010111011 : data_out = 24'b000000000011111101010100;
    16'b0000001010111100 : data_out = 24'b000000000011111101100100;
    16'b0000001010111101 : data_out = 24'b000000000011111101110100;
    16'b0000001010111110 : data_out = 24'b000000000011111110000011;
    16'b0000001010111111 : data_out = 24'b000000000011111110010011;
    16'b0000001011000000 : data_out = 24'b000000000011111110100011;
    16'b0000001011000001 : data_out = 24'b000000000011111110110011;
    16'b0000001011000010 : data_out = 24'b000000000011111111000011;
    16'b0000001011000011 : data_out = 24'b000000000011111111010011;
    16'b0000001011000100 : data_out = 24'b000000000011111111100011;
    16'b0000001011000101 : data_out = 24'b000000000011111111110011;
    16'b0000001011000110 : data_out = 24'b000000000100000000000011;
    16'b0000001011000111 : data_out = 24'b000000000100000000010011;
    16'b0000001011001000 : data_out = 24'b000000000100000000100011;
    16'b0000001011001001 : data_out = 24'b000000000100000000110011;
    16'b0000001011001010 : data_out = 24'b000000000100000001000011;
    16'b0000001011001011 : data_out = 24'b000000000100000001010011;
    16'b0000001011001100 : data_out = 24'b000000000100000001100011;
    16'b0000001011001101 : data_out = 24'b000000000100000001110011;
    16'b0000001011001110 : data_out = 24'b000000000100000010000100;
    16'b0000001011001111 : data_out = 24'b000000000100000010010100;
    16'b0000001011010000 : data_out = 24'b000000000100000010100100;
    16'b0000001011010001 : data_out = 24'b000000000100000010110100;
    16'b0000001011010010 : data_out = 24'b000000000100000011000100;
    16'b0000001011010011 : data_out = 24'b000000000100000011010100;
    16'b0000001011010100 : data_out = 24'b000000000100000011100101;
    16'b0000001011010101 : data_out = 24'b000000000100000011110101;
    16'b0000001011010110 : data_out = 24'b000000000100000100000101;
    16'b0000001011010111 : data_out = 24'b000000000100000100010101;
    16'b0000001011011000 : data_out = 24'b000000000100000100100110;
    16'b0000001011011001 : data_out = 24'b000000000100000100110110;
    16'b0000001011011010 : data_out = 24'b000000000100000101000110;
    16'b0000001011011011 : data_out = 24'b000000000100000101010111;
    16'b0000001011011100 : data_out = 24'b000000000100000101100111;
    16'b0000001011011101 : data_out = 24'b000000000100000101110111;
    16'b0000001011011110 : data_out = 24'b000000000100000110001000;
    16'b0000001011011111 : data_out = 24'b000000000100000110011000;
    16'b0000001011100000 : data_out = 24'b000000000100000110101000;
    16'b0000001011100001 : data_out = 24'b000000000100000110111001;
    16'b0000001011100010 : data_out = 24'b000000000100000111001001;
    16'b0000001011100011 : data_out = 24'b000000000100000111011010;
    16'b0000001011100100 : data_out = 24'b000000000100000111101010;
    16'b0000001011100101 : data_out = 24'b000000000100000111111011;
    16'b0000001011100110 : data_out = 24'b000000000100001000001011;
    16'b0000001011100111 : data_out = 24'b000000000100001000011100;
    16'b0000001011101000 : data_out = 24'b000000000100001000101100;
    16'b0000001011101001 : data_out = 24'b000000000100001000111101;
    16'b0000001011101010 : data_out = 24'b000000000100001001001101;
    16'b0000001011101011 : data_out = 24'b000000000100001001011110;
    16'b0000001011101100 : data_out = 24'b000000000100001001101111;
    16'b0000001011101101 : data_out = 24'b000000000100001001111111;
    16'b0000001011101110 : data_out = 24'b000000000100001010010000;
    16'b0000001011101111 : data_out = 24'b000000000100001010100000;
    16'b0000001011110000 : data_out = 24'b000000000100001010110001;
    16'b0000001011110001 : data_out = 24'b000000000100001011000010;
    16'b0000001011110010 : data_out = 24'b000000000100001011010010;
    16'b0000001011110011 : data_out = 24'b000000000100001011100011;
    16'b0000001011110100 : data_out = 24'b000000000100001011110100;
    16'b0000001011110101 : data_out = 24'b000000000100001100000101;
    16'b0000001011110110 : data_out = 24'b000000000100001100010101;
    16'b0000001011110111 : data_out = 24'b000000000100001100100110;
    16'b0000001011111000 : data_out = 24'b000000000100001100110111;
    16'b0000001011111001 : data_out = 24'b000000000100001101001000;
    16'b0000001011111010 : data_out = 24'b000000000100001101011001;
    16'b0000001011111011 : data_out = 24'b000000000100001101101001;
    16'b0000001011111100 : data_out = 24'b000000000100001101111010;
    16'b0000001011111101 : data_out = 24'b000000000100001110001011;
    16'b0000001011111110 : data_out = 24'b000000000100001110011100;
    16'b0000001011111111 : data_out = 24'b000000000100001110101101;
    16'b0000001100000000 : data_out = 24'b000000000100001110111110;
    16'b0000001100000001 : data_out = 24'b000000000100001111001111;
    16'b0000001100000010 : data_out = 24'b000000000100001111100000;
    16'b0000001100000011 : data_out = 24'b000000000100001111110001;
    16'b0000001100000100 : data_out = 24'b000000000100010000000010;
    16'b0000001100000101 : data_out = 24'b000000000100010000010011;
    16'b0000001100000110 : data_out = 24'b000000000100010000100100;
    16'b0000001100000111 : data_out = 24'b000000000100010000110101;
    16'b0000001100001000 : data_out = 24'b000000000100010001000110;
    16'b0000001100001001 : data_out = 24'b000000000100010001010111;
    16'b0000001100001010 : data_out = 24'b000000000100010001101000;
    16'b0000001100001011 : data_out = 24'b000000000100010001111001;
    16'b0000001100001100 : data_out = 24'b000000000100010010001010;
    16'b0000001100001101 : data_out = 24'b000000000100010010011100;
    16'b0000001100001110 : data_out = 24'b000000000100010010101101;
    16'b0000001100001111 : data_out = 24'b000000000100010010111110;
    16'b0000001100010000 : data_out = 24'b000000000100010011001111;
    16'b0000001100010001 : data_out = 24'b000000000100010011100000;
    16'b0000001100010010 : data_out = 24'b000000000100010011110010;
    16'b0000001100010011 : data_out = 24'b000000000100010100000011;
    16'b0000001100010100 : data_out = 24'b000000000100010100010100;
    16'b0000001100010101 : data_out = 24'b000000000100010100100101;
    16'b0000001100010110 : data_out = 24'b000000000100010100110111;
    16'b0000001100010111 : data_out = 24'b000000000100010101001000;
    16'b0000001100011000 : data_out = 24'b000000000100010101011001;
    16'b0000001100011001 : data_out = 24'b000000000100010101101011;
    16'b0000001100011010 : data_out = 24'b000000000100010101111100;
    16'b0000001100011011 : data_out = 24'b000000000100010110001101;
    16'b0000001100011100 : data_out = 24'b000000000100010110011111;
    16'b0000001100011101 : data_out = 24'b000000000100010110110000;
    16'b0000001100011110 : data_out = 24'b000000000100010111000010;
    16'b0000001100011111 : data_out = 24'b000000000100010111010011;
    16'b0000001100100000 : data_out = 24'b000000000100010111100100;
    16'b0000001100100001 : data_out = 24'b000000000100010111110110;
    16'b0000001100100010 : data_out = 24'b000000000100011000000111;
    16'b0000001100100011 : data_out = 24'b000000000100011000011001;
    16'b0000001100100100 : data_out = 24'b000000000100011000101011;
    16'b0000001100100101 : data_out = 24'b000000000100011000111100;
    16'b0000001100100110 : data_out = 24'b000000000100011001001110;
    16'b0000001100100111 : data_out = 24'b000000000100011001011111;
    16'b0000001100101000 : data_out = 24'b000000000100011001110001;
    16'b0000001100101001 : data_out = 24'b000000000100011010000010;
    16'b0000001100101010 : data_out = 24'b000000000100011010010100;
    16'b0000001100101011 : data_out = 24'b000000000100011010100110;
    16'b0000001100101100 : data_out = 24'b000000000100011010110111;
    16'b0000001100101101 : data_out = 24'b000000000100011011001001;
    16'b0000001100101110 : data_out = 24'b000000000100011011011011;
    16'b0000001100101111 : data_out = 24'b000000000100011011101101;
    16'b0000001100110000 : data_out = 24'b000000000100011011111110;
    16'b0000001100110001 : data_out = 24'b000000000100011100010000;
    16'b0000001100110010 : data_out = 24'b000000000100011100100010;
    16'b0000001100110011 : data_out = 24'b000000000100011100110100;
    16'b0000001100110100 : data_out = 24'b000000000100011101000101;
    16'b0000001100110101 : data_out = 24'b000000000100011101010111;
    16'b0000001100110110 : data_out = 24'b000000000100011101101001;
    16'b0000001100110111 : data_out = 24'b000000000100011101111011;
    16'b0000001100111000 : data_out = 24'b000000000100011110001101;
    16'b0000001100111001 : data_out = 24'b000000000100011110011111;
    16'b0000001100111010 : data_out = 24'b000000000100011110110001;
    16'b0000001100111011 : data_out = 24'b000000000100011111000011;
    16'b0000001100111100 : data_out = 24'b000000000100011111010100;
    16'b0000001100111101 : data_out = 24'b000000000100011111100110;
    16'b0000001100111110 : data_out = 24'b000000000100011111111000;
    16'b0000001100111111 : data_out = 24'b000000000100100000001010;
    16'b0000001101000000 : data_out = 24'b000000000100100000011100;
    16'b0000001101000001 : data_out = 24'b000000000100100000101110;
    16'b0000001101000010 : data_out = 24'b000000000100100001000001;
    16'b0000001101000011 : data_out = 24'b000000000100100001010011;
    16'b0000001101000100 : data_out = 24'b000000000100100001100101;
    16'b0000001101000101 : data_out = 24'b000000000100100001110111;
    16'b0000001101000110 : data_out = 24'b000000000100100010001001;
    16'b0000001101000111 : data_out = 24'b000000000100100010011011;
    16'b0000001101001000 : data_out = 24'b000000000100100010101101;
    16'b0000001101001001 : data_out = 24'b000000000100100010111111;
    16'b0000001101001010 : data_out = 24'b000000000100100011010010;
    16'b0000001101001011 : data_out = 24'b000000000100100011100100;
    16'b0000001101001100 : data_out = 24'b000000000100100011110110;
    16'b0000001101001101 : data_out = 24'b000000000100100100001000;
    16'b0000001101001110 : data_out = 24'b000000000100100100011011;
    16'b0000001101001111 : data_out = 24'b000000000100100100101101;
    16'b0000001101010000 : data_out = 24'b000000000100100100111111;
    16'b0000001101010001 : data_out = 24'b000000000100100101010001;
    16'b0000001101010010 : data_out = 24'b000000000100100101100100;
    16'b0000001101010011 : data_out = 24'b000000000100100101110110;
    16'b0000001101010100 : data_out = 24'b000000000100100110001001;
    16'b0000001101010101 : data_out = 24'b000000000100100110011011;
    16'b0000001101010110 : data_out = 24'b000000000100100110101101;
    16'b0000001101010111 : data_out = 24'b000000000100100111000000;
    16'b0000001101011000 : data_out = 24'b000000000100100111010010;
    16'b0000001101011001 : data_out = 24'b000000000100100111100101;
    16'b0000001101011010 : data_out = 24'b000000000100100111110111;
    16'b0000001101011011 : data_out = 24'b000000000100101000001010;
    16'b0000001101011100 : data_out = 24'b000000000100101000011100;
    16'b0000001101011101 : data_out = 24'b000000000100101000101111;
    16'b0000001101011110 : data_out = 24'b000000000100101001000001;
    16'b0000001101011111 : data_out = 24'b000000000100101001010100;
    16'b0000001101100000 : data_out = 24'b000000000100101001100110;
    16'b0000001101100001 : data_out = 24'b000000000100101001111001;
    16'b0000001101100010 : data_out = 24'b000000000100101010001100;
    16'b0000001101100011 : data_out = 24'b000000000100101010011110;
    16'b0000001101100100 : data_out = 24'b000000000100101010110001;
    16'b0000001101100101 : data_out = 24'b000000000100101011000100;
    16'b0000001101100110 : data_out = 24'b000000000100101011010110;
    16'b0000001101100111 : data_out = 24'b000000000100101011101001;
    16'b0000001101101000 : data_out = 24'b000000000100101011111100;
    16'b0000001101101001 : data_out = 24'b000000000100101100001111;
    16'b0000001101101010 : data_out = 24'b000000000100101100100001;
    16'b0000001101101011 : data_out = 24'b000000000100101100110100;
    16'b0000001101101100 : data_out = 24'b000000000100101101000111;
    16'b0000001101101101 : data_out = 24'b000000000100101101011010;
    16'b0000001101101110 : data_out = 24'b000000000100101101101101;
    16'b0000001101101111 : data_out = 24'b000000000100101110000000;
    16'b0000001101110000 : data_out = 24'b000000000100101110010010;
    16'b0000001101110001 : data_out = 24'b000000000100101110100101;
    16'b0000001101110010 : data_out = 24'b000000000100101110111000;
    16'b0000001101110011 : data_out = 24'b000000000100101111001011;
    16'b0000001101110100 : data_out = 24'b000000000100101111011110;
    16'b0000001101110101 : data_out = 24'b000000000100101111110001;
    16'b0000001101110110 : data_out = 24'b000000000100110000000100;
    16'b0000001101110111 : data_out = 24'b000000000100110000010111;
    16'b0000001101111000 : data_out = 24'b000000000100110000101010;
    16'b0000001101111001 : data_out = 24'b000000000100110000111101;
    16'b0000001101111010 : data_out = 24'b000000000100110001010000;
    16'b0000001101111011 : data_out = 24'b000000000100110001100011;
    16'b0000001101111100 : data_out = 24'b000000000100110001110110;
    16'b0000001101111101 : data_out = 24'b000000000100110010001010;
    16'b0000001101111110 : data_out = 24'b000000000100110010011101;
    16'b0000001101111111 : data_out = 24'b000000000100110010110000;
    16'b0000001110000000 : data_out = 24'b000000000100110011000011;
    16'b0000001110000001 : data_out = 24'b000000000100110011010110;
    16'b0000001110000010 : data_out = 24'b000000000100110011101010;
    16'b0000001110000011 : data_out = 24'b000000000100110011111101;
    16'b0000001110000100 : data_out = 24'b000000000100110100010000;
    16'b0000001110000101 : data_out = 24'b000000000100110100100011;
    16'b0000001110000110 : data_out = 24'b000000000100110100110111;
    16'b0000001110000111 : data_out = 24'b000000000100110101001010;
    16'b0000001110001000 : data_out = 24'b000000000100110101011101;
    16'b0000001110001001 : data_out = 24'b000000000100110101110001;
    16'b0000001110001010 : data_out = 24'b000000000100110110000100;
    16'b0000001110001011 : data_out = 24'b000000000100110110010111;
    16'b0000001110001100 : data_out = 24'b000000000100110110101011;
    16'b0000001110001101 : data_out = 24'b000000000100110110111110;
    16'b0000001110001110 : data_out = 24'b000000000100110111010010;
    16'b0000001110001111 : data_out = 24'b000000000100110111100101;
    16'b0000001110010000 : data_out = 24'b000000000100110111111001;
    16'b0000001110010001 : data_out = 24'b000000000100111000001100;
    16'b0000001110010010 : data_out = 24'b000000000100111000100000;
    16'b0000001110010011 : data_out = 24'b000000000100111000110011;
    16'b0000001110010100 : data_out = 24'b000000000100111001000111;
    16'b0000001110010101 : data_out = 24'b000000000100111001011010;
    16'b0000001110010110 : data_out = 24'b000000000100111001101110;
    16'b0000001110010111 : data_out = 24'b000000000100111010000001;
    16'b0000001110011000 : data_out = 24'b000000000100111010010101;
    16'b0000001110011001 : data_out = 24'b000000000100111010101001;
    16'b0000001110011010 : data_out = 24'b000000000100111010111100;
    16'b0000001110011011 : data_out = 24'b000000000100111011010000;
    16'b0000001110011100 : data_out = 24'b000000000100111011100100;
    16'b0000001110011101 : data_out = 24'b000000000100111011111000;
    16'b0000001110011110 : data_out = 24'b000000000100111100001011;
    16'b0000001110011111 : data_out = 24'b000000000100111100011111;
    16'b0000001110100000 : data_out = 24'b000000000100111100110011;
    16'b0000001110100001 : data_out = 24'b000000000100111101000111;
    16'b0000001110100010 : data_out = 24'b000000000100111101011011;
    16'b0000001110100011 : data_out = 24'b000000000100111101101110;
    16'b0000001110100100 : data_out = 24'b000000000100111110000010;
    16'b0000001110100101 : data_out = 24'b000000000100111110010110;
    16'b0000001110100110 : data_out = 24'b000000000100111110101010;
    16'b0000001110100111 : data_out = 24'b000000000100111110111110;
    16'b0000001110101000 : data_out = 24'b000000000100111111010010;
    16'b0000001110101001 : data_out = 24'b000000000100111111100110;
    16'b0000001110101010 : data_out = 24'b000000000100111111111010;
    16'b0000001110101011 : data_out = 24'b000000000101000000001110;
    16'b0000001110101100 : data_out = 24'b000000000101000000100010;
    16'b0000001110101101 : data_out = 24'b000000000101000000110110;
    16'b0000001110101110 : data_out = 24'b000000000101000001001010;
    16'b0000001110101111 : data_out = 24'b000000000101000001011110;
    16'b0000001110110000 : data_out = 24'b000000000101000001110010;
    16'b0000001110110001 : data_out = 24'b000000000101000010000110;
    16'b0000001110110010 : data_out = 24'b000000000101000010011010;
    16'b0000001110110011 : data_out = 24'b000000000101000010101111;
    16'b0000001110110100 : data_out = 24'b000000000101000011000011;
    16'b0000001110110101 : data_out = 24'b000000000101000011010111;
    16'b0000001110110110 : data_out = 24'b000000000101000011101011;
    16'b0000001110110111 : data_out = 24'b000000000101000011111111;
    16'b0000001110111000 : data_out = 24'b000000000101000100010100;
    16'b0000001110111001 : data_out = 24'b000000000101000100101000;
    16'b0000001110111010 : data_out = 24'b000000000101000100111100;
    16'b0000001110111011 : data_out = 24'b000000000101000101010001;
    16'b0000001110111100 : data_out = 24'b000000000101000101100101;
    16'b0000001110111101 : data_out = 24'b000000000101000101111001;
    16'b0000001110111110 : data_out = 24'b000000000101000110001110;
    16'b0000001110111111 : data_out = 24'b000000000101000110100010;
    16'b0000001111000000 : data_out = 24'b000000000101000110110111;
    16'b0000001111000001 : data_out = 24'b000000000101000111001011;
    16'b0000001111000010 : data_out = 24'b000000000101000111011111;
    16'b0000001111000011 : data_out = 24'b000000000101000111110100;
    16'b0000001111000100 : data_out = 24'b000000000101001000001000;
    16'b0000001111000101 : data_out = 24'b000000000101001000011101;
    16'b0000001111000110 : data_out = 24'b000000000101001000110001;
    16'b0000001111000111 : data_out = 24'b000000000101001001000110;
    16'b0000001111001000 : data_out = 24'b000000000101001001011011;
    16'b0000001111001001 : data_out = 24'b000000000101001001101111;
    16'b0000001111001010 : data_out = 24'b000000000101001010000100;
    16'b0000001111001011 : data_out = 24'b000000000101001010011000;
    16'b0000001111001100 : data_out = 24'b000000000101001010101101;
    16'b0000001111001101 : data_out = 24'b000000000101001011000010;
    16'b0000001111001110 : data_out = 24'b000000000101001011010110;
    16'b0000001111001111 : data_out = 24'b000000000101001011101011;
    16'b0000001111010000 : data_out = 24'b000000000101001100000000;
    16'b0000001111010001 : data_out = 24'b000000000101001100010101;
    16'b0000001111010010 : data_out = 24'b000000000101001100101001;
    16'b0000001111010011 : data_out = 24'b000000000101001100111110;
    16'b0000001111010100 : data_out = 24'b000000000101001101010011;
    16'b0000001111010101 : data_out = 24'b000000000101001101101000;
    16'b0000001111010110 : data_out = 24'b000000000101001101111101;
    16'b0000001111010111 : data_out = 24'b000000000101001110010010;
    16'b0000001111011000 : data_out = 24'b000000000101001110100111;
    16'b0000001111011001 : data_out = 24'b000000000101001110111100;
    16'b0000001111011010 : data_out = 24'b000000000101001111010000;
    16'b0000001111011011 : data_out = 24'b000000000101001111100101;
    16'b0000001111011100 : data_out = 24'b000000000101001111111010;
    16'b0000001111011101 : data_out = 24'b000000000101010000001111;
    16'b0000001111011110 : data_out = 24'b000000000101010000100100;
    16'b0000001111011111 : data_out = 24'b000000000101010000111001;
    16'b0000001111100000 : data_out = 24'b000000000101010001001111;
    16'b0000001111100001 : data_out = 24'b000000000101010001100100;
    16'b0000001111100010 : data_out = 24'b000000000101010001111001;
    16'b0000001111100011 : data_out = 24'b000000000101010010001110;
    16'b0000001111100100 : data_out = 24'b000000000101010010100011;
    16'b0000001111100101 : data_out = 24'b000000000101010010111000;
    16'b0000001111100110 : data_out = 24'b000000000101010011001101;
    16'b0000001111100111 : data_out = 24'b000000000101010011100011;
    16'b0000001111101000 : data_out = 24'b000000000101010011111000;
    16'b0000001111101001 : data_out = 24'b000000000101010100001101;
    16'b0000001111101010 : data_out = 24'b000000000101010100100010;
    16'b0000001111101011 : data_out = 24'b000000000101010100111000;
    16'b0000001111101100 : data_out = 24'b000000000101010101001101;
    16'b0000001111101101 : data_out = 24'b000000000101010101100010;
    16'b0000001111101110 : data_out = 24'b000000000101010101111000;
    16'b0000001111101111 : data_out = 24'b000000000101010110001101;
    16'b0000001111110000 : data_out = 24'b000000000101010110100010;
    16'b0000001111110001 : data_out = 24'b000000000101010110111000;
    16'b0000001111110010 : data_out = 24'b000000000101010111001101;
    16'b0000001111110011 : data_out = 24'b000000000101010111100011;
    16'b0000001111110100 : data_out = 24'b000000000101010111111000;
    16'b0000001111110101 : data_out = 24'b000000000101011000001110;
    16'b0000001111110110 : data_out = 24'b000000000101011000100011;
    16'b0000001111110111 : data_out = 24'b000000000101011000111001;
    16'b0000001111111000 : data_out = 24'b000000000101011001001110;
    16'b0000001111111001 : data_out = 24'b000000000101011001100100;
    16'b0000001111111010 : data_out = 24'b000000000101011001111010;
    16'b0000001111111011 : data_out = 24'b000000000101011010001111;
    16'b0000001111111100 : data_out = 24'b000000000101011010100101;
    16'b0000001111111101 : data_out = 24'b000000000101011010111011;
    16'b0000001111111110 : data_out = 24'b000000000101011011010000;
    16'b0000001111111111 : data_out = 24'b000000000101011011100110;
    16'b0000010000000000 : data_out = 24'b000000000101011011111100;
    16'b0000010000000001 : data_out = 24'b000000000101011100010001;
    16'b0000010000000010 : data_out = 24'b000000000101011100100111;
    16'b0000010000000011 : data_out = 24'b000000000101011100111101;
    16'b0000010000000100 : data_out = 24'b000000000101011101010011;
    16'b0000010000000101 : data_out = 24'b000000000101011101101001;
    16'b0000010000000110 : data_out = 24'b000000000101011101111111;
    16'b0000010000000111 : data_out = 24'b000000000101011110010100;
    16'b0000010000001000 : data_out = 24'b000000000101011110101010;
    16'b0000010000001001 : data_out = 24'b000000000101011111000000;
    16'b0000010000001010 : data_out = 24'b000000000101011111010110;
    16'b0000010000001011 : data_out = 24'b000000000101011111101100;
    16'b0000010000001100 : data_out = 24'b000000000101100000000010;
    16'b0000010000001101 : data_out = 24'b000000000101100000011000;
    16'b0000010000001110 : data_out = 24'b000000000101100000101110;
    16'b0000010000001111 : data_out = 24'b000000000101100001000100;
    16'b0000010000010000 : data_out = 24'b000000000101100001011010;
    16'b0000010000010001 : data_out = 24'b000000000101100001110000;
    16'b0000010000010010 : data_out = 24'b000000000101100010000111;
    16'b0000010000010011 : data_out = 24'b000000000101100010011101;
    16'b0000010000010100 : data_out = 24'b000000000101100010110011;
    16'b0000010000010101 : data_out = 24'b000000000101100011001001;
    16'b0000010000010110 : data_out = 24'b000000000101100011011111;
    16'b0000010000010111 : data_out = 24'b000000000101100011110101;
    16'b0000010000011000 : data_out = 24'b000000000101100100001100;
    16'b0000010000011001 : data_out = 24'b000000000101100100100010;
    16'b0000010000011010 : data_out = 24'b000000000101100100111000;
    16'b0000010000011011 : data_out = 24'b000000000101100101001111;
    16'b0000010000011100 : data_out = 24'b000000000101100101100101;
    16'b0000010000011101 : data_out = 24'b000000000101100101111011;
    16'b0000010000011110 : data_out = 24'b000000000101100110010010;
    16'b0000010000011111 : data_out = 24'b000000000101100110101000;
    16'b0000010000100000 : data_out = 24'b000000000101100110111111;
    16'b0000010000100001 : data_out = 24'b000000000101100111010101;
    16'b0000010000100010 : data_out = 24'b000000000101100111101011;
    16'b0000010000100011 : data_out = 24'b000000000101101000000010;
    16'b0000010000100100 : data_out = 24'b000000000101101000011000;
    16'b0000010000100101 : data_out = 24'b000000000101101000101111;
    16'b0000010000100110 : data_out = 24'b000000000101101001000110;
    16'b0000010000100111 : data_out = 24'b000000000101101001011100;
    16'b0000010000101000 : data_out = 24'b000000000101101001110011;
    16'b0000010000101001 : data_out = 24'b000000000101101010001001;
    16'b0000010000101010 : data_out = 24'b000000000101101010100000;
    16'b0000010000101011 : data_out = 24'b000000000101101010110111;
    16'b0000010000101100 : data_out = 24'b000000000101101011001101;
    16'b0000010000101101 : data_out = 24'b000000000101101011100100;
    16'b0000010000101110 : data_out = 24'b000000000101101011111011;
    16'b0000010000101111 : data_out = 24'b000000000101101100010010;
    16'b0000010000110000 : data_out = 24'b000000000101101100101000;
    16'b0000010000110001 : data_out = 24'b000000000101101100111111;
    16'b0000010000110010 : data_out = 24'b000000000101101101010110;
    16'b0000010000110011 : data_out = 24'b000000000101101101101101;
    16'b0000010000110100 : data_out = 24'b000000000101101110000100;
    16'b0000010000110101 : data_out = 24'b000000000101101110011011;
    16'b0000010000110110 : data_out = 24'b000000000101101110110001;
    16'b0000010000110111 : data_out = 24'b000000000101101111001000;
    16'b0000010000111000 : data_out = 24'b000000000101101111011111;
    16'b0000010000111001 : data_out = 24'b000000000101101111110110;
    16'b0000010000111010 : data_out = 24'b000000000101110000001101;
    16'b0000010000111011 : data_out = 24'b000000000101110000100100;
    16'b0000010000111100 : data_out = 24'b000000000101110000111011;
    16'b0000010000111101 : data_out = 24'b000000000101110001010010;
    16'b0000010000111110 : data_out = 24'b000000000101110001101010;
    16'b0000010000111111 : data_out = 24'b000000000101110010000001;
    16'b0000010001000000 : data_out = 24'b000000000101110010011000;
    16'b0000010001000001 : data_out = 24'b000000000101110010101111;
    16'b0000010001000010 : data_out = 24'b000000000101110011000110;
    16'b0000010001000011 : data_out = 24'b000000000101110011011101;
    16'b0000010001000100 : data_out = 24'b000000000101110011110101;
    16'b0000010001000101 : data_out = 24'b000000000101110100001100;
    16'b0000010001000110 : data_out = 24'b000000000101110100100011;
    16'b0000010001000111 : data_out = 24'b000000000101110100111010;
    16'b0000010001001000 : data_out = 24'b000000000101110101010010;
    16'b0000010001001001 : data_out = 24'b000000000101110101101001;
    16'b0000010001001010 : data_out = 24'b000000000101110110000000;
    16'b0000010001001011 : data_out = 24'b000000000101110110011000;
    16'b0000010001001100 : data_out = 24'b000000000101110110101111;
    16'b0000010001001101 : data_out = 24'b000000000101110111000111;
    16'b0000010001001110 : data_out = 24'b000000000101110111011110;
    16'b0000010001001111 : data_out = 24'b000000000101110111110110;
    16'b0000010001010000 : data_out = 24'b000000000101111000001101;
    16'b0000010001010001 : data_out = 24'b000000000101111000100101;
    16'b0000010001010010 : data_out = 24'b000000000101111000111100;
    16'b0000010001010011 : data_out = 24'b000000000101111001010100;
    16'b0000010001010100 : data_out = 24'b000000000101111001101011;
    16'b0000010001010101 : data_out = 24'b000000000101111010000011;
    16'b0000010001010110 : data_out = 24'b000000000101111010011011;
    16'b0000010001010111 : data_out = 24'b000000000101111010110010;
    16'b0000010001011000 : data_out = 24'b000000000101111011001010;
    16'b0000010001011001 : data_out = 24'b000000000101111011100010;
    16'b0000010001011010 : data_out = 24'b000000000101111011111001;
    16'b0000010001011011 : data_out = 24'b000000000101111100010001;
    16'b0000010001011100 : data_out = 24'b000000000101111100101001;
    16'b0000010001011101 : data_out = 24'b000000000101111101000001;
    16'b0000010001011110 : data_out = 24'b000000000101111101011001;
    16'b0000010001011111 : data_out = 24'b000000000101111101110000;
    16'b0000010001100000 : data_out = 24'b000000000101111110001000;
    16'b0000010001100001 : data_out = 24'b000000000101111110100000;
    16'b0000010001100010 : data_out = 24'b000000000101111110111000;
    16'b0000010001100011 : data_out = 24'b000000000101111111010000;
    16'b0000010001100100 : data_out = 24'b000000000101111111101000;
    16'b0000010001100101 : data_out = 24'b000000000110000000000000;
    16'b0000010001100110 : data_out = 24'b000000000110000000011000;
    16'b0000010001100111 : data_out = 24'b000000000110000000110000;
    16'b0000010001101000 : data_out = 24'b000000000110000001001000;
    16'b0000010001101001 : data_out = 24'b000000000110000001100000;
    16'b0000010001101010 : data_out = 24'b000000000110000001111000;
    16'b0000010001101011 : data_out = 24'b000000000110000010010000;
    16'b0000010001101100 : data_out = 24'b000000000110000010101001;
    16'b0000010001101101 : data_out = 24'b000000000110000011000001;
    16'b0000010001101110 : data_out = 24'b000000000110000011011001;
    16'b0000010001101111 : data_out = 24'b000000000110000011110001;
    16'b0000010001110000 : data_out = 24'b000000000110000100001001;
    16'b0000010001110001 : data_out = 24'b000000000110000100100010;
    16'b0000010001110010 : data_out = 24'b000000000110000100111010;
    16'b0000010001110011 : data_out = 24'b000000000110000101010010;
    16'b0000010001110100 : data_out = 24'b000000000110000101101011;
    16'b0000010001110101 : data_out = 24'b000000000110000110000011;
    16'b0000010001110110 : data_out = 24'b000000000110000110011011;
    16'b0000010001110111 : data_out = 24'b000000000110000110110100;
    16'b0000010001111000 : data_out = 24'b000000000110000111001100;
    16'b0000010001111001 : data_out = 24'b000000000110000111100101;
    16'b0000010001111010 : data_out = 24'b000000000110000111111101;
    16'b0000010001111011 : data_out = 24'b000000000110001000010110;
    16'b0000010001111100 : data_out = 24'b000000000110001000101110;
    16'b0000010001111101 : data_out = 24'b000000000110001001000111;
    16'b0000010001111110 : data_out = 24'b000000000110001001011111;
    16'b0000010001111111 : data_out = 24'b000000000110001001111000;
    16'b0000010010000000 : data_out = 24'b000000000110001010010001;
    16'b0000010010000001 : data_out = 24'b000000000110001010101001;
    16'b0000010010000010 : data_out = 24'b000000000110001011000010;
    16'b0000010010000011 : data_out = 24'b000000000110001011011011;
    16'b0000010010000100 : data_out = 24'b000000000110001011110011;
    16'b0000010010000101 : data_out = 24'b000000000110001100001100;
    16'b0000010010000110 : data_out = 24'b000000000110001100100101;
    16'b0000010010000111 : data_out = 24'b000000000110001100111110;
    16'b0000010010001000 : data_out = 24'b000000000110001101010111;
    16'b0000010010001001 : data_out = 24'b000000000110001101101111;
    16'b0000010010001010 : data_out = 24'b000000000110001110001000;
    16'b0000010010001011 : data_out = 24'b000000000110001110100001;
    16'b0000010010001100 : data_out = 24'b000000000110001110111010;
    16'b0000010010001101 : data_out = 24'b000000000110001111010011;
    16'b0000010010001110 : data_out = 24'b000000000110001111101100;
    16'b0000010010001111 : data_out = 24'b000000000110010000000101;
    16'b0000010010010000 : data_out = 24'b000000000110010000011110;
    16'b0000010010010001 : data_out = 24'b000000000110010000110111;
    16'b0000010010010010 : data_out = 24'b000000000110010001010000;
    16'b0000010010010011 : data_out = 24'b000000000110010001101001;
    16'b0000010010010100 : data_out = 24'b000000000110010010000010;
    16'b0000010010010101 : data_out = 24'b000000000110010010011011;
    16'b0000010010010110 : data_out = 24'b000000000110010010110101;
    16'b0000010010010111 : data_out = 24'b000000000110010011001110;
    16'b0000010010011000 : data_out = 24'b000000000110010011100111;
    16'b0000010010011001 : data_out = 24'b000000000110010100000000;
    16'b0000010010011010 : data_out = 24'b000000000110010100011010;
    16'b0000010010011011 : data_out = 24'b000000000110010100110011;
    16'b0000010010011100 : data_out = 24'b000000000110010101001100;
    16'b0000010010011101 : data_out = 24'b000000000110010101100101;
    16'b0000010010011110 : data_out = 24'b000000000110010101111111;
    16'b0000010010011111 : data_out = 24'b000000000110010110011000;
    16'b0000010010100000 : data_out = 24'b000000000110010110110010;
    16'b0000010010100001 : data_out = 24'b000000000110010111001011;
    16'b0000010010100010 : data_out = 24'b000000000110010111100101;
    16'b0000010010100011 : data_out = 24'b000000000110010111111110;
    16'b0000010010100100 : data_out = 24'b000000000110011000011000;
    16'b0000010010100101 : data_out = 24'b000000000110011000110001;
    16'b0000010010100110 : data_out = 24'b000000000110011001001011;
    16'b0000010010100111 : data_out = 24'b000000000110011001100100;
    16'b0000010010101000 : data_out = 24'b000000000110011001111110;
    16'b0000010010101001 : data_out = 24'b000000000110011010010111;
    16'b0000010010101010 : data_out = 24'b000000000110011010110001;
    16'b0000010010101011 : data_out = 24'b000000000110011011001011;
    16'b0000010010101100 : data_out = 24'b000000000110011011100101;
    16'b0000010010101101 : data_out = 24'b000000000110011011111110;
    16'b0000010010101110 : data_out = 24'b000000000110011100011000;
    16'b0000010010101111 : data_out = 24'b000000000110011100110010;
    16'b0000010010110000 : data_out = 24'b000000000110011101001100;
    16'b0000010010110001 : data_out = 24'b000000000110011101100101;
    16'b0000010010110010 : data_out = 24'b000000000110011101111111;
    16'b0000010010110011 : data_out = 24'b000000000110011110011001;
    16'b0000010010110100 : data_out = 24'b000000000110011110110011;
    16'b0000010010110101 : data_out = 24'b000000000110011111001101;
    16'b0000010010110110 : data_out = 24'b000000000110011111100111;
    16'b0000010010110111 : data_out = 24'b000000000110100000000001;
    16'b0000010010111000 : data_out = 24'b000000000110100000011011;
    16'b0000010010111001 : data_out = 24'b000000000110100000110101;
    16'b0000010010111010 : data_out = 24'b000000000110100001001111;
    16'b0000010010111011 : data_out = 24'b000000000110100001101001;
    16'b0000010010111100 : data_out = 24'b000000000110100010000011;
    16'b0000010010111101 : data_out = 24'b000000000110100010011101;
    16'b0000010010111110 : data_out = 24'b000000000110100010111000;
    16'b0000010010111111 : data_out = 24'b000000000110100011010010;
    16'b0000010011000000 : data_out = 24'b000000000110100011101100;
    16'b0000010011000001 : data_out = 24'b000000000110100100000110;
    16'b0000010011000010 : data_out = 24'b000000000110100100100001;
    16'b0000010011000011 : data_out = 24'b000000000110100100111011;
    16'b0000010011000100 : data_out = 24'b000000000110100101010101;
    16'b0000010011000101 : data_out = 24'b000000000110100101110000;
    16'b0000010011000110 : data_out = 24'b000000000110100110001010;
    16'b0000010011000111 : data_out = 24'b000000000110100110100100;
    16'b0000010011001000 : data_out = 24'b000000000110100110111111;
    16'b0000010011001001 : data_out = 24'b000000000110100111011001;
    16'b0000010011001010 : data_out = 24'b000000000110100111110100;
    16'b0000010011001011 : data_out = 24'b000000000110101000001110;
    16'b0000010011001100 : data_out = 24'b000000000110101000101001;
    16'b0000010011001101 : data_out = 24'b000000000110101001000011;
    16'b0000010011001110 : data_out = 24'b000000000110101001011110;
    16'b0000010011001111 : data_out = 24'b000000000110101001111000;
    16'b0000010011010000 : data_out = 24'b000000000110101010010011;
    16'b0000010011010001 : data_out = 24'b000000000110101010101110;
    16'b0000010011010010 : data_out = 24'b000000000110101011001000;
    16'b0000010011010011 : data_out = 24'b000000000110101011100011;
    16'b0000010011010100 : data_out = 24'b000000000110101011111110;
    16'b0000010011010101 : data_out = 24'b000000000110101100011001;
    16'b0000010011010110 : data_out = 24'b000000000110101100110011;
    16'b0000010011010111 : data_out = 24'b000000000110101101001110;
    16'b0000010011011000 : data_out = 24'b000000000110101101101001;
    16'b0000010011011001 : data_out = 24'b000000000110101110000100;
    16'b0000010011011010 : data_out = 24'b000000000110101110011111;
    16'b0000010011011011 : data_out = 24'b000000000110101110111010;
    16'b0000010011011100 : data_out = 24'b000000000110101111010101;
    16'b0000010011011101 : data_out = 24'b000000000110101111110000;
    16'b0000010011011110 : data_out = 24'b000000000110110000001011;
    16'b0000010011011111 : data_out = 24'b000000000110110000100110;
    16'b0000010011100000 : data_out = 24'b000000000110110001000001;
    16'b0000010011100001 : data_out = 24'b000000000110110001011100;
    16'b0000010011100010 : data_out = 24'b000000000110110001110111;
    16'b0000010011100011 : data_out = 24'b000000000110110010010010;
    16'b0000010011100100 : data_out = 24'b000000000110110010101101;
    16'b0000010011100101 : data_out = 24'b000000000110110011001000;
    16'b0000010011100110 : data_out = 24'b000000000110110011100100;
    16'b0000010011100111 : data_out = 24'b000000000110110011111111;
    16'b0000010011101000 : data_out = 24'b000000000110110100011010;
    16'b0000010011101001 : data_out = 24'b000000000110110100110101;
    16'b0000010011101010 : data_out = 24'b000000000110110101010001;
    16'b0000010011101011 : data_out = 24'b000000000110110101101100;
    16'b0000010011101100 : data_out = 24'b000000000110110110000111;
    16'b0000010011101101 : data_out = 24'b000000000110110110100011;
    16'b0000010011101110 : data_out = 24'b000000000110110110111110;
    16'b0000010011101111 : data_out = 24'b000000000110110111011010;
    16'b0000010011110000 : data_out = 24'b000000000110110111110101;
    16'b0000010011110001 : data_out = 24'b000000000110111000010001;
    16'b0000010011110010 : data_out = 24'b000000000110111000101100;
    16'b0000010011110011 : data_out = 24'b000000000110111001001000;
    16'b0000010011110100 : data_out = 24'b000000000110111001100011;
    16'b0000010011110101 : data_out = 24'b000000000110111001111111;
    16'b0000010011110110 : data_out = 24'b000000000110111010011011;
    16'b0000010011110111 : data_out = 24'b000000000110111010110110;
    16'b0000010011111000 : data_out = 24'b000000000110111011010010;
    16'b0000010011111001 : data_out = 24'b000000000110111011101110;
    16'b0000010011111010 : data_out = 24'b000000000110111100001001;
    16'b0000010011111011 : data_out = 24'b000000000110111100100101;
    16'b0000010011111100 : data_out = 24'b000000000110111101000001;
    16'b0000010011111101 : data_out = 24'b000000000110111101011101;
    16'b0000010011111110 : data_out = 24'b000000000110111101111001;
    16'b0000010011111111 : data_out = 24'b000000000110111110010100;
    16'b0000010100000000 : data_out = 24'b000000000110111110110000;
    16'b0000010100000001 : data_out = 24'b000000000110111111001100;
    16'b0000010100000010 : data_out = 24'b000000000110111111101000;
    16'b0000010100000011 : data_out = 24'b000000000111000000000100;
    16'b0000010100000100 : data_out = 24'b000000000111000000100000;
    16'b0000010100000101 : data_out = 24'b000000000111000000111100;
    16'b0000010100000110 : data_out = 24'b000000000111000001011000;
    16'b0000010100000111 : data_out = 24'b000000000111000001110101;
    16'b0000010100001000 : data_out = 24'b000000000111000010010001;
    16'b0000010100001001 : data_out = 24'b000000000111000010101101;
    16'b0000010100001010 : data_out = 24'b000000000111000011001001;
    16'b0000010100001011 : data_out = 24'b000000000111000011100101;
    16'b0000010100001100 : data_out = 24'b000000000111000100000001;
    16'b0000010100001101 : data_out = 24'b000000000111000100011110;
    16'b0000010100001110 : data_out = 24'b000000000111000100111010;
    16'b0000010100001111 : data_out = 24'b000000000111000101010110;
    16'b0000010100010000 : data_out = 24'b000000000111000101110011;
    16'b0000010100010001 : data_out = 24'b000000000111000110001111;
    16'b0000010100010010 : data_out = 24'b000000000111000110101011;
    16'b0000010100010011 : data_out = 24'b000000000111000111001000;
    16'b0000010100010100 : data_out = 24'b000000000111000111100100;
    16'b0000010100010101 : data_out = 24'b000000000111001000000001;
    16'b0000010100010110 : data_out = 24'b000000000111001000011101;
    16'b0000010100010111 : data_out = 24'b000000000111001000111010;
    16'b0000010100011000 : data_out = 24'b000000000111001001010110;
    16'b0000010100011001 : data_out = 24'b000000000111001001110011;
    16'b0000010100011010 : data_out = 24'b000000000111001010010000;
    16'b0000010100011011 : data_out = 24'b000000000111001010101100;
    16'b0000010100011100 : data_out = 24'b000000000111001011001001;
    16'b0000010100011101 : data_out = 24'b000000000111001011100110;
    16'b0000010100011110 : data_out = 24'b000000000111001100000010;
    16'b0000010100011111 : data_out = 24'b000000000111001100011111;
    16'b0000010100100000 : data_out = 24'b000000000111001100111100;
    16'b0000010100100001 : data_out = 24'b000000000111001101011001;
    16'b0000010100100010 : data_out = 24'b000000000111001101110110;
    16'b0000010100100011 : data_out = 24'b000000000111001110010011;
    16'b0000010100100100 : data_out = 24'b000000000111001110101111;
    16'b0000010100100101 : data_out = 24'b000000000111001111001100;
    16'b0000010100100110 : data_out = 24'b000000000111001111101001;
    16'b0000010100100111 : data_out = 24'b000000000111010000000110;
    16'b0000010100101000 : data_out = 24'b000000000111010000100011;
    16'b0000010100101001 : data_out = 24'b000000000111010001000000;
    16'b0000010100101010 : data_out = 24'b000000000111010001011110;
    16'b0000010100101011 : data_out = 24'b000000000111010001111011;
    16'b0000010100101100 : data_out = 24'b000000000111010010011000;
    16'b0000010100101101 : data_out = 24'b000000000111010010110101;
    16'b0000010100101110 : data_out = 24'b000000000111010011010010;
    16'b0000010100101111 : data_out = 24'b000000000111010011101111;
    16'b0000010100110000 : data_out = 24'b000000000111010100001101;
    16'b0000010100110001 : data_out = 24'b000000000111010100101010;
    16'b0000010100110010 : data_out = 24'b000000000111010101000111;
    16'b0000010100110011 : data_out = 24'b000000000111010101100101;
    16'b0000010100110100 : data_out = 24'b000000000111010110000010;
    16'b0000010100110101 : data_out = 24'b000000000111010110011111;
    16'b0000010100110110 : data_out = 24'b000000000111010110111101;
    16'b0000010100110111 : data_out = 24'b000000000111010111011010;
    16'b0000010100111000 : data_out = 24'b000000000111010111111000;
    16'b0000010100111001 : data_out = 24'b000000000111011000010101;
    16'b0000010100111010 : data_out = 24'b000000000111011000110011;
    16'b0000010100111011 : data_out = 24'b000000000111011001010000;
    16'b0000010100111100 : data_out = 24'b000000000111011001101110;
    16'b0000010100111101 : data_out = 24'b000000000111011010001011;
    16'b0000010100111110 : data_out = 24'b000000000111011010101001;
    16'b0000010100111111 : data_out = 24'b000000000111011011000111;
    16'b0000010101000000 : data_out = 24'b000000000111011011100100;
    16'b0000010101000001 : data_out = 24'b000000000111011100000010;
    16'b0000010101000010 : data_out = 24'b000000000111011100100000;
    16'b0000010101000011 : data_out = 24'b000000000111011100111110;
    16'b0000010101000100 : data_out = 24'b000000000111011101011100;
    16'b0000010101000101 : data_out = 24'b000000000111011101111001;
    16'b0000010101000110 : data_out = 24'b000000000111011110010111;
    16'b0000010101000111 : data_out = 24'b000000000111011110110101;
    16'b0000010101001000 : data_out = 24'b000000000111011111010011;
    16'b0000010101001001 : data_out = 24'b000000000111011111110001;
    16'b0000010101001010 : data_out = 24'b000000000111100000001111;
    16'b0000010101001011 : data_out = 24'b000000000111100000101101;
    16'b0000010101001100 : data_out = 24'b000000000111100001001011;
    16'b0000010101001101 : data_out = 24'b000000000111100001101001;
    16'b0000010101001110 : data_out = 24'b000000000111100010000111;
    16'b0000010101001111 : data_out = 24'b000000000111100010100110;
    16'b0000010101010000 : data_out = 24'b000000000111100011000100;
    16'b0000010101010001 : data_out = 24'b000000000111100011100010;
    16'b0000010101010010 : data_out = 24'b000000000111100100000000;
    16'b0000010101010011 : data_out = 24'b000000000111100100011110;
    16'b0000010101010100 : data_out = 24'b000000000111100100111101;
    16'b0000010101010101 : data_out = 24'b000000000111100101011011;
    16'b0000010101010110 : data_out = 24'b000000000111100101111001;
    16'b0000010101010111 : data_out = 24'b000000000111100110011000;
    16'b0000010101011000 : data_out = 24'b000000000111100110110110;
    16'b0000010101011001 : data_out = 24'b000000000111100111010101;
    16'b0000010101011010 : data_out = 24'b000000000111100111110011;
    16'b0000010101011011 : data_out = 24'b000000000111101000010010;
    16'b0000010101011100 : data_out = 24'b000000000111101000110000;
    16'b0000010101011101 : data_out = 24'b000000000111101001001111;
    16'b0000010101011110 : data_out = 24'b000000000111101001101101;
    16'b0000010101011111 : data_out = 24'b000000000111101010001100;
    16'b0000010101100000 : data_out = 24'b000000000111101010101011;
    16'b0000010101100001 : data_out = 24'b000000000111101011001001;
    16'b0000010101100010 : data_out = 24'b000000000111101011101000;
    16'b0000010101100011 : data_out = 24'b000000000111101100000111;
    16'b0000010101100100 : data_out = 24'b000000000111101100100110;
    16'b0000010101100101 : data_out = 24'b000000000111101101000100;
    16'b0000010101100110 : data_out = 24'b000000000111101101100011;
    16'b0000010101100111 : data_out = 24'b000000000111101110000010;
    16'b0000010101101000 : data_out = 24'b000000000111101110100001;
    16'b0000010101101001 : data_out = 24'b000000000111101111000000;
    16'b0000010101101010 : data_out = 24'b000000000111101111011111;
    16'b0000010101101011 : data_out = 24'b000000000111101111111110;
    16'b0000010101101100 : data_out = 24'b000000000111110000011101;
    16'b0000010101101101 : data_out = 24'b000000000111110000111100;
    16'b0000010101101110 : data_out = 24'b000000000111110001011011;
    16'b0000010101101111 : data_out = 24'b000000000111110001111010;
    16'b0000010101110000 : data_out = 24'b000000000111110010011001;
    16'b0000010101110001 : data_out = 24'b000000000111110010111000;
    16'b0000010101110010 : data_out = 24'b000000000111110011011000;
    16'b0000010101110011 : data_out = 24'b000000000111110011110111;
    16'b0000010101110100 : data_out = 24'b000000000111110100010110;
    16'b0000010101110101 : data_out = 24'b000000000111110100110101;
    16'b0000010101110110 : data_out = 24'b000000000111110101010101;
    16'b0000010101110111 : data_out = 24'b000000000111110101110100;
    16'b0000010101111000 : data_out = 24'b000000000111110110010011;
    16'b0000010101111001 : data_out = 24'b000000000111110110110011;
    16'b0000010101111010 : data_out = 24'b000000000111110111010010;
    16'b0000010101111011 : data_out = 24'b000000000111110111110010;
    16'b0000010101111100 : data_out = 24'b000000000111111000010001;
    16'b0000010101111101 : data_out = 24'b000000000111111000110001;
    16'b0000010101111110 : data_out = 24'b000000000111111001010000;
    16'b0000010101111111 : data_out = 24'b000000000111111001110000;
    16'b0000010110000000 : data_out = 24'b000000000111111010001111;
    16'b0000010110000001 : data_out = 24'b000000000111111010101111;
    16'b0000010110000010 : data_out = 24'b000000000111111011001111;
    16'b0000010110000011 : data_out = 24'b000000000111111011101111;
    16'b0000010110000100 : data_out = 24'b000000000111111100001110;
    16'b0000010110000101 : data_out = 24'b000000000111111100101110;
    16'b0000010110000110 : data_out = 24'b000000000111111101001110;
    16'b0000010110000111 : data_out = 24'b000000000111111101101110;
    16'b0000010110001000 : data_out = 24'b000000000111111110001110;
    16'b0000010110001001 : data_out = 24'b000000000111111110101110;
    16'b0000010110001010 : data_out = 24'b000000000111111111001101;
    16'b0000010110001011 : data_out = 24'b000000000111111111101101;
    16'b0000010110001100 : data_out = 24'b000000001000000000001101;
    16'b0000010110001101 : data_out = 24'b000000001000000000101101;
    16'b0000010110001110 : data_out = 24'b000000001000000001001101;
    16'b0000010110001111 : data_out = 24'b000000001000000001101110;
    16'b0000010110010000 : data_out = 24'b000000001000000010001110;
    16'b0000010110010001 : data_out = 24'b000000001000000010101110;
    16'b0000010110010010 : data_out = 24'b000000001000000011001110;
    16'b0000010110010011 : data_out = 24'b000000001000000011101110;
    16'b0000010110010100 : data_out = 24'b000000001000000100001111;
    16'b0000010110010101 : data_out = 24'b000000001000000100101111;
    16'b0000010110010110 : data_out = 24'b000000001000000101001111;
    16'b0000010110010111 : data_out = 24'b000000001000000101101111;
    16'b0000010110011000 : data_out = 24'b000000001000000110010000;
    16'b0000010110011001 : data_out = 24'b000000001000000110110000;
    16'b0000010110011010 : data_out = 24'b000000001000000111010001;
    16'b0000010110011011 : data_out = 24'b000000001000000111110001;
    16'b0000010110011100 : data_out = 24'b000000001000001000010010;
    16'b0000010110011101 : data_out = 24'b000000001000001000110010;
    16'b0000010110011110 : data_out = 24'b000000001000001001010011;
    16'b0000010110011111 : data_out = 24'b000000001000001001110011;
    16'b0000010110100000 : data_out = 24'b000000001000001010010100;
    16'b0000010110100001 : data_out = 24'b000000001000001010110101;
    16'b0000010110100010 : data_out = 24'b000000001000001011010101;
    16'b0000010110100011 : data_out = 24'b000000001000001011110110;
    16'b0000010110100100 : data_out = 24'b000000001000001100010111;
    16'b0000010110100101 : data_out = 24'b000000001000001100111000;
    16'b0000010110100110 : data_out = 24'b000000001000001101011000;
    16'b0000010110100111 : data_out = 24'b000000001000001101111001;
    16'b0000010110101000 : data_out = 24'b000000001000001110011010;
    16'b0000010110101001 : data_out = 24'b000000001000001110111011;
    16'b0000010110101010 : data_out = 24'b000000001000001111011100;
    16'b0000010110101011 : data_out = 24'b000000001000001111111101;
    16'b0000010110101100 : data_out = 24'b000000001000010000011110;
    16'b0000010110101101 : data_out = 24'b000000001000010000111111;
    16'b0000010110101110 : data_out = 24'b000000001000010001100000;
    16'b0000010110101111 : data_out = 24'b000000001000010010000001;
    16'b0000010110110000 : data_out = 24'b000000001000010010100010;
    16'b0000010110110001 : data_out = 24'b000000001000010011000100;
    16'b0000010110110010 : data_out = 24'b000000001000010011100101;
    16'b0000010110110011 : data_out = 24'b000000001000010100000110;
    16'b0000010110110100 : data_out = 24'b000000001000010100100111;
    16'b0000010110110101 : data_out = 24'b000000001000010101001001;
    16'b0000010110110110 : data_out = 24'b000000001000010101101010;
    16'b0000010110110111 : data_out = 24'b000000001000010110001011;
    16'b0000010110111000 : data_out = 24'b000000001000010110101101;
    16'b0000010110111001 : data_out = 24'b000000001000010111001110;
    16'b0000010110111010 : data_out = 24'b000000001000010111110000;
    16'b0000010110111011 : data_out = 24'b000000001000011000010001;
    16'b0000010110111100 : data_out = 24'b000000001000011000110011;
    16'b0000010110111101 : data_out = 24'b000000001000011001010100;
    16'b0000010110111110 : data_out = 24'b000000001000011001110110;
    16'b0000010110111111 : data_out = 24'b000000001000011010010111;
    16'b0000010111000000 : data_out = 24'b000000001000011010111001;
    16'b0000010111000001 : data_out = 24'b000000001000011011011011;
    16'b0000010111000010 : data_out = 24'b000000001000011011111101;
    16'b0000010111000011 : data_out = 24'b000000001000011100011110;
    16'b0000010111000100 : data_out = 24'b000000001000011101000000;
    16'b0000010111000101 : data_out = 24'b000000001000011101100010;
    16'b0000010111000110 : data_out = 24'b000000001000011110000100;
    16'b0000010111000111 : data_out = 24'b000000001000011110100110;
    16'b0000010111001000 : data_out = 24'b000000001000011111001000;
    16'b0000010111001001 : data_out = 24'b000000001000011111101010;
    16'b0000010111001010 : data_out = 24'b000000001000100000001100;
    16'b0000010111001011 : data_out = 24'b000000001000100000101110;
    16'b0000010111001100 : data_out = 24'b000000001000100001010000;
    16'b0000010111001101 : data_out = 24'b000000001000100001110010;
    16'b0000010111001110 : data_out = 24'b000000001000100010010100;
    16'b0000010111001111 : data_out = 24'b000000001000100010110110;
    16'b0000010111010000 : data_out = 24'b000000001000100011011000;
    16'b0000010111010001 : data_out = 24'b000000001000100011111010;
    16'b0000010111010010 : data_out = 24'b000000001000100100011101;
    16'b0000010111010011 : data_out = 24'b000000001000100100111111;
    16'b0000010111010100 : data_out = 24'b000000001000100101100001;
    16'b0000010111010101 : data_out = 24'b000000001000100110000100;
    16'b0000010111010110 : data_out = 24'b000000001000100110100110;
    16'b0000010111010111 : data_out = 24'b000000001000100111001001;
    16'b0000010111011000 : data_out = 24'b000000001000100111101011;
    16'b0000010111011001 : data_out = 24'b000000001000101000001110;
    16'b0000010111011010 : data_out = 24'b000000001000101000110000;
    16'b0000010111011011 : data_out = 24'b000000001000101001010011;
    16'b0000010111011100 : data_out = 24'b000000001000101001110101;
    16'b0000010111011101 : data_out = 24'b000000001000101010011000;
    16'b0000010111011110 : data_out = 24'b000000001000101010111010;
    16'b0000010111011111 : data_out = 24'b000000001000101011011101;
    16'b0000010111100000 : data_out = 24'b000000001000101100000000;
    16'b0000010111100001 : data_out = 24'b000000001000101100100011;
    16'b0000010111100010 : data_out = 24'b000000001000101101000101;
    16'b0000010111100011 : data_out = 24'b000000001000101101101000;
    16'b0000010111100100 : data_out = 24'b000000001000101110001011;
    16'b0000010111100101 : data_out = 24'b000000001000101110101110;
    16'b0000010111100110 : data_out = 24'b000000001000101111010001;
    16'b0000010111100111 : data_out = 24'b000000001000101111110100;
    16'b0000010111101000 : data_out = 24'b000000001000110000010111;
    16'b0000010111101001 : data_out = 24'b000000001000110000111010;
    16'b0000010111101010 : data_out = 24'b000000001000110001011101;
    16'b0000010111101011 : data_out = 24'b000000001000110010000000;
    16'b0000010111101100 : data_out = 24'b000000001000110010100011;
    16'b0000010111101101 : data_out = 24'b000000001000110011000111;
    16'b0000010111101110 : data_out = 24'b000000001000110011101010;
    16'b0000010111101111 : data_out = 24'b000000001000110100001101;
    16'b0000010111110000 : data_out = 24'b000000001000110100110000;
    16'b0000010111110001 : data_out = 24'b000000001000110101010100;
    16'b0000010111110010 : data_out = 24'b000000001000110101110111;
    16'b0000010111110011 : data_out = 24'b000000001000110110011010;
    16'b0000010111110100 : data_out = 24'b000000001000110110111110;
    16'b0000010111110101 : data_out = 24'b000000001000110111100001;
    16'b0000010111110110 : data_out = 24'b000000001000111000000101;
    16'b0000010111110111 : data_out = 24'b000000001000111000101000;
    16'b0000010111111000 : data_out = 24'b000000001000111001001100;
    16'b0000010111111001 : data_out = 24'b000000001000111001101111;
    16'b0000010111111010 : data_out = 24'b000000001000111010010011;
    16'b0000010111111011 : data_out = 24'b000000001000111010110111;
    16'b0000010111111100 : data_out = 24'b000000001000111011011010;
    16'b0000010111111101 : data_out = 24'b000000001000111011111110;
    16'b0000010111111110 : data_out = 24'b000000001000111100100010;
    16'b0000010111111111 : data_out = 24'b000000001000111101000110;
    16'b0000011000000000 : data_out = 24'b000000001000111101101001;
    16'b0000011000000001 : data_out = 24'b000000001000111110001101;
    16'b0000011000000010 : data_out = 24'b000000001000111110110001;
    16'b0000011000000011 : data_out = 24'b000000001000111111010101;
    16'b0000011000000100 : data_out = 24'b000000001000111111111001;
    16'b0000011000000101 : data_out = 24'b000000001001000000011101;
    16'b0000011000000110 : data_out = 24'b000000001001000001000001;
    16'b0000011000000111 : data_out = 24'b000000001001000001100101;
    16'b0000011000001000 : data_out = 24'b000000001001000010001001;
    16'b0000011000001001 : data_out = 24'b000000001001000010101110;
    16'b0000011000001010 : data_out = 24'b000000001001000011010010;
    16'b0000011000001011 : data_out = 24'b000000001001000011110110;
    16'b0000011000001100 : data_out = 24'b000000001001000100011010;
    16'b0000011000001101 : data_out = 24'b000000001001000100111111;
    16'b0000011000001110 : data_out = 24'b000000001001000101100011;
    16'b0000011000001111 : data_out = 24'b000000001001000110000111;
    16'b0000011000010000 : data_out = 24'b000000001001000110101100;
    16'b0000011000010001 : data_out = 24'b000000001001000111010000;
    16'b0000011000010010 : data_out = 24'b000000001001000111110101;
    16'b0000011000010011 : data_out = 24'b000000001001001000011001;
    16'b0000011000010100 : data_out = 24'b000000001001001000111110;
    16'b0000011000010101 : data_out = 24'b000000001001001001100010;
    16'b0000011000010110 : data_out = 24'b000000001001001010000111;
    16'b0000011000010111 : data_out = 24'b000000001001001010101011;
    16'b0000011000011000 : data_out = 24'b000000001001001011010000;
    16'b0000011000011001 : data_out = 24'b000000001001001011110101;
    16'b0000011000011010 : data_out = 24'b000000001001001100011010;
    16'b0000011000011011 : data_out = 24'b000000001001001100111110;
    16'b0000011000011100 : data_out = 24'b000000001001001101100011;
    16'b0000011000011101 : data_out = 24'b000000001001001110001000;
    16'b0000011000011110 : data_out = 24'b000000001001001110101101;
    16'b0000011000011111 : data_out = 24'b000000001001001111010010;
    16'b0000011000100000 : data_out = 24'b000000001001001111110111;
    16'b0000011000100001 : data_out = 24'b000000001001010000011100;
    16'b0000011000100010 : data_out = 24'b000000001001010001000001;
    16'b0000011000100011 : data_out = 24'b000000001001010001100110;
    16'b0000011000100100 : data_out = 24'b000000001001010010001011;
    16'b0000011000100101 : data_out = 24'b000000001001010010110000;
    16'b0000011000100110 : data_out = 24'b000000001001010011010110;
    16'b0000011000100111 : data_out = 24'b000000001001010011111011;
    16'b0000011000101000 : data_out = 24'b000000001001010100100000;
    16'b0000011000101001 : data_out = 24'b000000001001010101000101;
    16'b0000011000101010 : data_out = 24'b000000001001010101101011;
    16'b0000011000101011 : data_out = 24'b000000001001010110010000;
    16'b0000011000101100 : data_out = 24'b000000001001010110110101;
    16'b0000011000101101 : data_out = 24'b000000001001010111011011;
    16'b0000011000101110 : data_out = 24'b000000001001011000000000;
    16'b0000011000101111 : data_out = 24'b000000001001011000100110;
    16'b0000011000110000 : data_out = 24'b000000001001011001001011;
    16'b0000011000110001 : data_out = 24'b000000001001011001110001;
    16'b0000011000110010 : data_out = 24'b000000001001011010010111;
    16'b0000011000110011 : data_out = 24'b000000001001011010111100;
    16'b0000011000110100 : data_out = 24'b000000001001011011100010;
    16'b0000011000110101 : data_out = 24'b000000001001011100001000;
    16'b0000011000110110 : data_out = 24'b000000001001011100101110;
    16'b0000011000110111 : data_out = 24'b000000001001011101010011;
    16'b0000011000111000 : data_out = 24'b000000001001011101111001;
    16'b0000011000111001 : data_out = 24'b000000001001011110011111;
    16'b0000011000111010 : data_out = 24'b000000001001011111000101;
    16'b0000011000111011 : data_out = 24'b000000001001011111101011;
    16'b0000011000111100 : data_out = 24'b000000001001100000010001;
    16'b0000011000111101 : data_out = 24'b000000001001100000110111;
    16'b0000011000111110 : data_out = 24'b000000001001100001011101;
    16'b0000011000111111 : data_out = 24'b000000001001100010000011;
    16'b0000011001000000 : data_out = 24'b000000001001100010101001;
    16'b0000011001000001 : data_out = 24'b000000001001100011010000;
    16'b0000011001000010 : data_out = 24'b000000001001100011110110;
    16'b0000011001000011 : data_out = 24'b000000001001100100011100;
    16'b0000011001000100 : data_out = 24'b000000001001100101000010;
    16'b0000011001000101 : data_out = 24'b000000001001100101101001;
    16'b0000011001000110 : data_out = 24'b000000001001100110001111;
    16'b0000011001000111 : data_out = 24'b000000001001100110110101;
    16'b0000011001001000 : data_out = 24'b000000001001100111011100;
    16'b0000011001001001 : data_out = 24'b000000001001101000000010;
    16'b0000011001001010 : data_out = 24'b000000001001101000101001;
    16'b0000011001001011 : data_out = 24'b000000001001101001001111;
    16'b0000011001001100 : data_out = 24'b000000001001101001110110;
    16'b0000011001001101 : data_out = 24'b000000001001101010011101;
    16'b0000011001001110 : data_out = 24'b000000001001101011000011;
    16'b0000011001001111 : data_out = 24'b000000001001101011101010;
    16'b0000011001010000 : data_out = 24'b000000001001101100010001;
    16'b0000011001010001 : data_out = 24'b000000001001101100111000;
    16'b0000011001010010 : data_out = 24'b000000001001101101011110;
    16'b0000011001010011 : data_out = 24'b000000001001101110000101;
    16'b0000011001010100 : data_out = 24'b000000001001101110101100;
    16'b0000011001010101 : data_out = 24'b000000001001101111010011;
    16'b0000011001010110 : data_out = 24'b000000001001101111111010;
    16'b0000011001010111 : data_out = 24'b000000001001110000100001;
    16'b0000011001011000 : data_out = 24'b000000001001110001001000;
    16'b0000011001011001 : data_out = 24'b000000001001110001101111;
    16'b0000011001011010 : data_out = 24'b000000001001110010010110;
    16'b0000011001011011 : data_out = 24'b000000001001110010111110;
    16'b0000011001011100 : data_out = 24'b000000001001110011100101;
    16'b0000011001011101 : data_out = 24'b000000001001110100001100;
    16'b0000011001011110 : data_out = 24'b000000001001110100110011;
    16'b0000011001011111 : data_out = 24'b000000001001110101011011;
    16'b0000011001100000 : data_out = 24'b000000001001110110000010;
    16'b0000011001100001 : data_out = 24'b000000001001110110101001;
    16'b0000011001100010 : data_out = 24'b000000001001110111010001;
    16'b0000011001100011 : data_out = 24'b000000001001110111111000;
    16'b0000011001100100 : data_out = 24'b000000001001111000100000;
    16'b0000011001100101 : data_out = 24'b000000001001111001000111;
    16'b0000011001100110 : data_out = 24'b000000001001111001101111;
    16'b0000011001100111 : data_out = 24'b000000001001111010010111;
    16'b0000011001101000 : data_out = 24'b000000001001111010111110;
    16'b0000011001101001 : data_out = 24'b000000001001111011100110;
    16'b0000011001101010 : data_out = 24'b000000001001111100001110;
    16'b0000011001101011 : data_out = 24'b000000001001111100110101;
    16'b0000011001101100 : data_out = 24'b000000001001111101011101;
    16'b0000011001101101 : data_out = 24'b000000001001111110000101;
    16'b0000011001101110 : data_out = 24'b000000001001111110101101;
    16'b0000011001101111 : data_out = 24'b000000001001111111010101;
    16'b0000011001110000 : data_out = 24'b000000001001111111111101;
    16'b0000011001110001 : data_out = 24'b000000001010000000100101;
    16'b0000011001110010 : data_out = 24'b000000001010000001001101;
    16'b0000011001110011 : data_out = 24'b000000001010000001110101;
    16'b0000011001110100 : data_out = 24'b000000001010000010011101;
    16'b0000011001110101 : data_out = 24'b000000001010000011000101;
    16'b0000011001110110 : data_out = 24'b000000001010000011101110;
    16'b0000011001110111 : data_out = 24'b000000001010000100010110;
    16'b0000011001111000 : data_out = 24'b000000001010000100111110;
    16'b0000011001111001 : data_out = 24'b000000001010000101100110;
    16'b0000011001111010 : data_out = 24'b000000001010000110001111;
    16'b0000011001111011 : data_out = 24'b000000001010000110110111;
    16'b0000011001111100 : data_out = 24'b000000001010000111100000;
    16'b0000011001111101 : data_out = 24'b000000001010001000001000;
    16'b0000011001111110 : data_out = 24'b000000001010001000110001;
    16'b0000011001111111 : data_out = 24'b000000001010001001011001;
    16'b0000011010000000 : data_out = 24'b000000001010001010000010;
    16'b0000011010000001 : data_out = 24'b000000001010001010101011;
    16'b0000011010000010 : data_out = 24'b000000001010001011010011;
    16'b0000011010000011 : data_out = 24'b000000001010001011111100;
    16'b0000011010000100 : data_out = 24'b000000001010001100100101;
    16'b0000011010000101 : data_out = 24'b000000001010001101001110;
    16'b0000011010000110 : data_out = 24'b000000001010001101110110;
    16'b0000011010000111 : data_out = 24'b000000001010001110011111;
    16'b0000011010001000 : data_out = 24'b000000001010001111001000;
    16'b0000011010001001 : data_out = 24'b000000001010001111110001;
    16'b0000011010001010 : data_out = 24'b000000001010010000011010;
    16'b0000011010001011 : data_out = 24'b000000001010010001000011;
    16'b0000011010001100 : data_out = 24'b000000001010010001101100;
    16'b0000011010001101 : data_out = 24'b000000001010010010010101;
    16'b0000011010001110 : data_out = 24'b000000001010010010111111;
    16'b0000011010001111 : data_out = 24'b000000001010010011101000;
    16'b0000011010010000 : data_out = 24'b000000001010010100010001;
    16'b0000011010010001 : data_out = 24'b000000001010010100111010;
    16'b0000011010010010 : data_out = 24'b000000001010010101100100;
    16'b0000011010010011 : data_out = 24'b000000001010010110001101;
    16'b0000011010010100 : data_out = 24'b000000001010010110110110;
    16'b0000011010010101 : data_out = 24'b000000001010010111100000;
    16'b0000011010010110 : data_out = 24'b000000001010011000001001;
    16'b0000011010010111 : data_out = 24'b000000001010011000110011;
    16'b0000011010011000 : data_out = 24'b000000001010011001011100;
    16'b0000011010011001 : data_out = 24'b000000001010011010000110;
    16'b0000011010011010 : data_out = 24'b000000001010011010110000;
    16'b0000011010011011 : data_out = 24'b000000001010011011011001;
    16'b0000011010011100 : data_out = 24'b000000001010011100000011;
    16'b0000011010011101 : data_out = 24'b000000001010011100101101;
    16'b0000011010011110 : data_out = 24'b000000001010011101010111;
    16'b0000011010011111 : data_out = 24'b000000001010011110000001;
    16'b0000011010100000 : data_out = 24'b000000001010011110101011;
    16'b0000011010100001 : data_out = 24'b000000001010011111010100;
    16'b0000011010100010 : data_out = 24'b000000001010011111111110;
    16'b0000011010100011 : data_out = 24'b000000001010100000101000;
    16'b0000011010100100 : data_out = 24'b000000001010100001010011;
    16'b0000011010100101 : data_out = 24'b000000001010100001111101;
    16'b0000011010100110 : data_out = 24'b000000001010100010100111;
    16'b0000011010100111 : data_out = 24'b000000001010100011010001;
    16'b0000011010101000 : data_out = 24'b000000001010100011111011;
    16'b0000011010101001 : data_out = 24'b000000001010100100100101;
    16'b0000011010101010 : data_out = 24'b000000001010100101010000;
    16'b0000011010101011 : data_out = 24'b000000001010100101111010;
    16'b0000011010101100 : data_out = 24'b000000001010100110100100;
    16'b0000011010101101 : data_out = 24'b000000001010100111001111;
    16'b0000011010101110 : data_out = 24'b000000001010100111111001;
    16'b0000011010101111 : data_out = 24'b000000001010101000100100;
    16'b0000011010110000 : data_out = 24'b000000001010101001001110;
    16'b0000011010110001 : data_out = 24'b000000001010101001111001;
    16'b0000011010110010 : data_out = 24'b000000001010101010100100;
    16'b0000011010110011 : data_out = 24'b000000001010101011001110;
    16'b0000011010110100 : data_out = 24'b000000001010101011111001;
    16'b0000011010110101 : data_out = 24'b000000001010101100100100;
    16'b0000011010110110 : data_out = 24'b000000001010101101001111;
    16'b0000011010110111 : data_out = 24'b000000001010101101111010;
    16'b0000011010111000 : data_out = 24'b000000001010101110100100;
    16'b0000011010111001 : data_out = 24'b000000001010101111001111;
    16'b0000011010111010 : data_out = 24'b000000001010101111111010;
    16'b0000011010111011 : data_out = 24'b000000001010110000100101;
    16'b0000011010111100 : data_out = 24'b000000001010110001010000;
    16'b0000011010111101 : data_out = 24'b000000001010110001111011;
    16'b0000011010111110 : data_out = 24'b000000001010110010100111;
    16'b0000011010111111 : data_out = 24'b000000001010110011010010;
    16'b0000011011000000 : data_out = 24'b000000001010110011111101;
    16'b0000011011000001 : data_out = 24'b000000001010110100101000;
    16'b0000011011000010 : data_out = 24'b000000001010110101010100;
    16'b0000011011000011 : data_out = 24'b000000001010110101111111;
    16'b0000011011000100 : data_out = 24'b000000001010110110101010;
    16'b0000011011000101 : data_out = 24'b000000001010110111010110;
    16'b0000011011000110 : data_out = 24'b000000001010111000000001;
    16'b0000011011000111 : data_out = 24'b000000001010111000101101;
    16'b0000011011001000 : data_out = 24'b000000001010111001011000;
    16'b0000011011001001 : data_out = 24'b000000001010111010000100;
    16'b0000011011001010 : data_out = 24'b000000001010111010110000;
    16'b0000011011001011 : data_out = 24'b000000001010111011011011;
    16'b0000011011001100 : data_out = 24'b000000001010111100000111;
    16'b0000011011001101 : data_out = 24'b000000001010111100110011;
    16'b0000011011001110 : data_out = 24'b000000001010111101011111;
    16'b0000011011001111 : data_out = 24'b000000001010111110001011;
    16'b0000011011010000 : data_out = 24'b000000001010111110110110;
    16'b0000011011010001 : data_out = 24'b000000001010111111100010;
    16'b0000011011010010 : data_out = 24'b000000001011000000001110;
    16'b0000011011010011 : data_out = 24'b000000001011000000111010;
    16'b0000011011010100 : data_out = 24'b000000001011000001100110;
    16'b0000011011010101 : data_out = 24'b000000001011000010010011;
    16'b0000011011010110 : data_out = 24'b000000001011000010111111;
    16'b0000011011010111 : data_out = 24'b000000001011000011101011;
    16'b0000011011011000 : data_out = 24'b000000001011000100010111;
    16'b0000011011011001 : data_out = 24'b000000001011000101000100;
    16'b0000011011011010 : data_out = 24'b000000001011000101110000;
    16'b0000011011011011 : data_out = 24'b000000001011000110011100;
    16'b0000011011011100 : data_out = 24'b000000001011000111001001;
    16'b0000011011011101 : data_out = 24'b000000001011000111110101;
    16'b0000011011011110 : data_out = 24'b000000001011001000100010;
    16'b0000011011011111 : data_out = 24'b000000001011001001001110;
    16'b0000011011100000 : data_out = 24'b000000001011001001111011;
    16'b0000011011100001 : data_out = 24'b000000001011001010100111;
    16'b0000011011100010 : data_out = 24'b000000001011001011010100;
    16'b0000011011100011 : data_out = 24'b000000001011001100000001;
    16'b0000011011100100 : data_out = 24'b000000001011001100101110;
    16'b0000011011100101 : data_out = 24'b000000001011001101011010;
    16'b0000011011100110 : data_out = 24'b000000001011001110000111;
    16'b0000011011100111 : data_out = 24'b000000001011001110110100;
    16'b0000011011101000 : data_out = 24'b000000001011001111100001;
    16'b0000011011101001 : data_out = 24'b000000001011010000001110;
    16'b0000011011101010 : data_out = 24'b000000001011010000111011;
    16'b0000011011101011 : data_out = 24'b000000001011010001101000;
    16'b0000011011101100 : data_out = 24'b000000001011010010010101;
    16'b0000011011101101 : data_out = 24'b000000001011010011000011;
    16'b0000011011101110 : data_out = 24'b000000001011010011110000;
    16'b0000011011101111 : data_out = 24'b000000001011010100011101;
    16'b0000011011110000 : data_out = 24'b000000001011010101001010;
    16'b0000011011110001 : data_out = 24'b000000001011010101111000;
    16'b0000011011110010 : data_out = 24'b000000001011010110100101;
    16'b0000011011110011 : data_out = 24'b000000001011010111010011;
    16'b0000011011110100 : data_out = 24'b000000001011011000000000;
    16'b0000011011110101 : data_out = 24'b000000001011011000101110;
    16'b0000011011110110 : data_out = 24'b000000001011011001011011;
    16'b0000011011110111 : data_out = 24'b000000001011011010001001;
    16'b0000011011111000 : data_out = 24'b000000001011011010110110;
    16'b0000011011111001 : data_out = 24'b000000001011011011100100;
    16'b0000011011111010 : data_out = 24'b000000001011011100010010;
    16'b0000011011111011 : data_out = 24'b000000001011011101000000;
    16'b0000011011111100 : data_out = 24'b000000001011011101101101;
    16'b0000011011111101 : data_out = 24'b000000001011011110011011;
    16'b0000011011111110 : data_out = 24'b000000001011011111001001;
    16'b0000011011111111 : data_out = 24'b000000001011011111110111;
    16'b0000011100000000 : data_out = 24'b000000001011100000100101;
    16'b0000011100000001 : data_out = 24'b000000001011100001010011;
    16'b0000011100000010 : data_out = 24'b000000001011100010000001;
    16'b0000011100000011 : data_out = 24'b000000001011100010110000;
    16'b0000011100000100 : data_out = 24'b000000001011100011011110;
    16'b0000011100000101 : data_out = 24'b000000001011100100001100;
    16'b0000011100000110 : data_out = 24'b000000001011100100111010;
    16'b0000011100000111 : data_out = 24'b000000001011100101101001;
    16'b0000011100001000 : data_out = 24'b000000001011100110010111;
    16'b0000011100001001 : data_out = 24'b000000001011100111000101;
    16'b0000011100001010 : data_out = 24'b000000001011100111110100;
    16'b0000011100001011 : data_out = 24'b000000001011101000100010;
    16'b0000011100001100 : data_out = 24'b000000001011101001010001;
    16'b0000011100001101 : data_out = 24'b000000001011101001111111;
    16'b0000011100001110 : data_out = 24'b000000001011101010101110;
    16'b0000011100001111 : data_out = 24'b000000001011101011011101;
    16'b0000011100010000 : data_out = 24'b000000001011101100001100;
    16'b0000011100010001 : data_out = 24'b000000001011101100111010;
    16'b0000011100010010 : data_out = 24'b000000001011101101101001;
    16'b0000011100010011 : data_out = 24'b000000001011101110011000;
    16'b0000011100010100 : data_out = 24'b000000001011101111000111;
    16'b0000011100010101 : data_out = 24'b000000001011101111110110;
    16'b0000011100010110 : data_out = 24'b000000001011110000100101;
    16'b0000011100010111 : data_out = 24'b000000001011110001010100;
    16'b0000011100011000 : data_out = 24'b000000001011110010000011;
    16'b0000011100011001 : data_out = 24'b000000001011110010110010;
    16'b0000011100011010 : data_out = 24'b000000001011110011100001;
    16'b0000011100011011 : data_out = 24'b000000001011110100010001;
    16'b0000011100011100 : data_out = 24'b000000001011110101000000;
    16'b0000011100011101 : data_out = 24'b000000001011110101101111;
    16'b0000011100011110 : data_out = 24'b000000001011110110011111;
    16'b0000011100011111 : data_out = 24'b000000001011110111001110;
    16'b0000011100100000 : data_out = 24'b000000001011110111111110;
    16'b0000011100100001 : data_out = 24'b000000001011111000101101;
    16'b0000011100100010 : data_out = 24'b000000001011111001011101;
    16'b0000011100100011 : data_out = 24'b000000001011111010001100;
    16'b0000011100100100 : data_out = 24'b000000001011111010111100;
    16'b0000011100100101 : data_out = 24'b000000001011111011101100;
    16'b0000011100100110 : data_out = 24'b000000001011111100011011;
    16'b0000011100100111 : data_out = 24'b000000001011111101001011;
    16'b0000011100101000 : data_out = 24'b000000001011111101111011;
    16'b0000011100101001 : data_out = 24'b000000001011111110101011;
    16'b0000011100101010 : data_out = 24'b000000001011111111011011;
    16'b0000011100101011 : data_out = 24'b000000001100000000001011;
    16'b0000011100101100 : data_out = 24'b000000001100000000111011;
    16'b0000011100101101 : data_out = 24'b000000001100000001101011;
    16'b0000011100101110 : data_out = 24'b000000001100000010011011;
    16'b0000011100101111 : data_out = 24'b000000001100000011001011;
    16'b0000011100110000 : data_out = 24'b000000001100000011111100;
    16'b0000011100110001 : data_out = 24'b000000001100000100101100;
    16'b0000011100110010 : data_out = 24'b000000001100000101011100;
    16'b0000011100110011 : data_out = 24'b000000001100000110001101;
    16'b0000011100110100 : data_out = 24'b000000001100000110111101;
    16'b0000011100110101 : data_out = 24'b000000001100000111101101;
    16'b0000011100110110 : data_out = 24'b000000001100001000011110;
    16'b0000011100110111 : data_out = 24'b000000001100001001001110;
    16'b0000011100111000 : data_out = 24'b000000001100001001111111;
    16'b0000011100111001 : data_out = 24'b000000001100001010110000;
    16'b0000011100111010 : data_out = 24'b000000001100001011100000;
    16'b0000011100111011 : data_out = 24'b000000001100001100010001;
    16'b0000011100111100 : data_out = 24'b000000001100001101000010;
    16'b0000011100111101 : data_out = 24'b000000001100001101110011;
    16'b0000011100111110 : data_out = 24'b000000001100001110100100;
    16'b0000011100111111 : data_out = 24'b000000001100001111010101;
    16'b0000011101000000 : data_out = 24'b000000001100010000000110;
    16'b0000011101000001 : data_out = 24'b000000001100010000110111;
    16'b0000011101000010 : data_out = 24'b000000001100010001101000;
    16'b0000011101000011 : data_out = 24'b000000001100010010011001;
    16'b0000011101000100 : data_out = 24'b000000001100010011001010;
    16'b0000011101000101 : data_out = 24'b000000001100010011111011;
    16'b0000011101000110 : data_out = 24'b000000001100010100101100;
    16'b0000011101000111 : data_out = 24'b000000001100010101011110;
    16'b0000011101001000 : data_out = 24'b000000001100010110001111;
    16'b0000011101001001 : data_out = 24'b000000001100010111000001;
    16'b0000011101001010 : data_out = 24'b000000001100010111110010;
    16'b0000011101001011 : data_out = 24'b000000001100011000100100;
    16'b0000011101001100 : data_out = 24'b000000001100011001010101;
    16'b0000011101001101 : data_out = 24'b000000001100011010000111;
    16'b0000011101001110 : data_out = 24'b000000001100011010111000;
    16'b0000011101001111 : data_out = 24'b000000001100011011101010;
    16'b0000011101010000 : data_out = 24'b000000001100011100011100;
    16'b0000011101010001 : data_out = 24'b000000001100011101001110;
    16'b0000011101010010 : data_out = 24'b000000001100011101111111;
    16'b0000011101010011 : data_out = 24'b000000001100011110110001;
    16'b0000011101010100 : data_out = 24'b000000001100011111100011;
    16'b0000011101010101 : data_out = 24'b000000001100100000010101;
    16'b0000011101010110 : data_out = 24'b000000001100100001000111;
    16'b0000011101010111 : data_out = 24'b000000001100100001111001;
    16'b0000011101011000 : data_out = 24'b000000001100100010101100;
    16'b0000011101011001 : data_out = 24'b000000001100100011011110;
    16'b0000011101011010 : data_out = 24'b000000001100100100010000;
    16'b0000011101011011 : data_out = 24'b000000001100100101000010;
    16'b0000011101011100 : data_out = 24'b000000001100100101110101;
    16'b0000011101011101 : data_out = 24'b000000001100100110100111;
    16'b0000011101011110 : data_out = 24'b000000001100100111011010;
    16'b0000011101011111 : data_out = 24'b000000001100101000001100;
    16'b0000011101100000 : data_out = 24'b000000001100101000111111;
    16'b0000011101100001 : data_out = 24'b000000001100101001110001;
    16'b0000011101100010 : data_out = 24'b000000001100101010100100;
    16'b0000011101100011 : data_out = 24'b000000001100101011010110;
    16'b0000011101100100 : data_out = 24'b000000001100101100001001;
    16'b0000011101100101 : data_out = 24'b000000001100101100111100;
    16'b0000011101100110 : data_out = 24'b000000001100101101101111;
    16'b0000011101100111 : data_out = 24'b000000001100101110100010;
    16'b0000011101101000 : data_out = 24'b000000001100101111010101;
    16'b0000011101101001 : data_out = 24'b000000001100110000001000;
    16'b0000011101101010 : data_out = 24'b000000001100110000111011;
    16'b0000011101101011 : data_out = 24'b000000001100110001101110;
    16'b0000011101101100 : data_out = 24'b000000001100110010100001;
    16'b0000011101101101 : data_out = 24'b000000001100110011010100;
    16'b0000011101101110 : data_out = 24'b000000001100110100000111;
    16'b0000011101101111 : data_out = 24'b000000001100110100111011;
    16'b0000011101110000 : data_out = 24'b000000001100110101101110;
    16'b0000011101110001 : data_out = 24'b000000001100110110100001;
    16'b0000011101110010 : data_out = 24'b000000001100110111010101;
    16'b0000011101110011 : data_out = 24'b000000001100111000001000;
    16'b0000011101110100 : data_out = 24'b000000001100111000111100;
    16'b0000011101110101 : data_out = 24'b000000001100111001101111;
    16'b0000011101110110 : data_out = 24'b000000001100111010100011;
    16'b0000011101110111 : data_out = 24'b000000001100111011010111;
    16'b0000011101111000 : data_out = 24'b000000001100111100001010;
    16'b0000011101111001 : data_out = 24'b000000001100111100111110;
    16'b0000011101111010 : data_out = 24'b000000001100111101110010;
    16'b0000011101111011 : data_out = 24'b000000001100111110100110;
    16'b0000011101111100 : data_out = 24'b000000001100111111011010;
    16'b0000011101111101 : data_out = 24'b000000001101000000001110;
    16'b0000011101111110 : data_out = 24'b000000001101000001000010;
    16'b0000011101111111 : data_out = 24'b000000001101000001110110;
    16'b0000011110000000 : data_out = 24'b000000001101000010101010;
    16'b0000011110000001 : data_out = 24'b000000001101000011011110;
    16'b0000011110000010 : data_out = 24'b000000001101000100010010;
    16'b0000011110000011 : data_out = 24'b000000001101000101000111;
    16'b0000011110000100 : data_out = 24'b000000001101000101111011;
    16'b0000011110000101 : data_out = 24'b000000001101000110110000;
    16'b0000011110000110 : data_out = 24'b000000001101000111100100;
    16'b0000011110000111 : data_out = 24'b000000001101001000011000;
    16'b0000011110001000 : data_out = 24'b000000001101001001001101;
    16'b0000011110001001 : data_out = 24'b000000001101001010000010;
    16'b0000011110001010 : data_out = 24'b000000001101001010110110;
    16'b0000011110001011 : data_out = 24'b000000001101001011101011;
    16'b0000011110001100 : data_out = 24'b000000001101001100100000;
    16'b0000011110001101 : data_out = 24'b000000001101001101010101;
    16'b0000011110001110 : data_out = 24'b000000001101001110001001;
    16'b0000011110001111 : data_out = 24'b000000001101001110111110;
    16'b0000011110010000 : data_out = 24'b000000001101001111110011;
    16'b0000011110010001 : data_out = 24'b000000001101010000101000;
    16'b0000011110010010 : data_out = 24'b000000001101010001011101;
    16'b0000011110010011 : data_out = 24'b000000001101010010010010;
    16'b0000011110010100 : data_out = 24'b000000001101010011001000;
    16'b0000011110010101 : data_out = 24'b000000001101010011111101;
    16'b0000011110010110 : data_out = 24'b000000001101010100110010;
    16'b0000011110010111 : data_out = 24'b000000001101010101100111;
    16'b0000011110011000 : data_out = 24'b000000001101010110011101;
    16'b0000011110011001 : data_out = 24'b000000001101010111010010;
    16'b0000011110011010 : data_out = 24'b000000001101011000001000;
    16'b0000011110011011 : data_out = 24'b000000001101011000111101;
    16'b0000011110011100 : data_out = 24'b000000001101011001110011;
    16'b0000011110011101 : data_out = 24'b000000001101011010101001;
    16'b0000011110011110 : data_out = 24'b000000001101011011011110;
    16'b0000011110011111 : data_out = 24'b000000001101011100010100;
    16'b0000011110100000 : data_out = 24'b000000001101011101001010;
    16'b0000011110100001 : data_out = 24'b000000001101011110000000;
    16'b0000011110100010 : data_out = 24'b000000001101011110110101;
    16'b0000011110100011 : data_out = 24'b000000001101011111101011;
    16'b0000011110100100 : data_out = 24'b000000001101100000100001;
    16'b0000011110100101 : data_out = 24'b000000001101100001011000;
    16'b0000011110100110 : data_out = 24'b000000001101100010001110;
    16'b0000011110100111 : data_out = 24'b000000001101100011000100;
    16'b0000011110101000 : data_out = 24'b000000001101100011111010;
    16'b0000011110101001 : data_out = 24'b000000001101100100110000;
    16'b0000011110101010 : data_out = 24'b000000001101100101100111;
    16'b0000011110101011 : data_out = 24'b000000001101100110011101;
    16'b0000011110101100 : data_out = 24'b000000001101100111010011;
    16'b0000011110101101 : data_out = 24'b000000001101101000001010;
    16'b0000011110101110 : data_out = 24'b000000001101101001000000;
    16'b0000011110101111 : data_out = 24'b000000001101101001110111;
    16'b0000011110110000 : data_out = 24'b000000001101101010101110;
    16'b0000011110110001 : data_out = 24'b000000001101101011100100;
    16'b0000011110110010 : data_out = 24'b000000001101101100011011;
    16'b0000011110110011 : data_out = 24'b000000001101101101010010;
    16'b0000011110110100 : data_out = 24'b000000001101101110001001;
    16'b0000011110110101 : data_out = 24'b000000001101101111000000;
    16'b0000011110110110 : data_out = 24'b000000001101101111110111;
    16'b0000011110110111 : data_out = 24'b000000001101110000101110;
    16'b0000011110111000 : data_out = 24'b000000001101110001100101;
    16'b0000011110111001 : data_out = 24'b000000001101110010011100;
    16'b0000011110111010 : data_out = 24'b000000001101110011010011;
    16'b0000011110111011 : data_out = 24'b000000001101110100001010;
    16'b0000011110111100 : data_out = 24'b000000001101110101000010;
    16'b0000011110111101 : data_out = 24'b000000001101110101111001;
    16'b0000011110111110 : data_out = 24'b000000001101110110110000;
    16'b0000011110111111 : data_out = 24'b000000001101110111101000;
    16'b0000011111000000 : data_out = 24'b000000001101111000011111;
    16'b0000011111000001 : data_out = 24'b000000001101111001010111;
    16'b0000011111000010 : data_out = 24'b000000001101111010001110;
    16'b0000011111000011 : data_out = 24'b000000001101111011000110;
    16'b0000011111000100 : data_out = 24'b000000001101111011111110;
    16'b0000011111000101 : data_out = 24'b000000001101111100110110;
    16'b0000011111000110 : data_out = 24'b000000001101111101101101;
    16'b0000011111000111 : data_out = 24'b000000001101111110100101;
    16'b0000011111001000 : data_out = 24'b000000001101111111011101;
    16'b0000011111001001 : data_out = 24'b000000001110000000010101;
    16'b0000011111001010 : data_out = 24'b000000001110000001001101;
    16'b0000011111001011 : data_out = 24'b000000001110000010000101;
    16'b0000011111001100 : data_out = 24'b000000001110000010111110;
    16'b0000011111001101 : data_out = 24'b000000001110000011110110;
    16'b0000011111001110 : data_out = 24'b000000001110000100101110;
    16'b0000011111001111 : data_out = 24'b000000001110000101100110;
    16'b0000011111010000 : data_out = 24'b000000001110000110011111;
    16'b0000011111010001 : data_out = 24'b000000001110000111010111;
    16'b0000011111010010 : data_out = 24'b000000001110001000010000;
    16'b0000011111010011 : data_out = 24'b000000001110001001001000;
    16'b0000011111010100 : data_out = 24'b000000001110001010000001;
    16'b0000011111010101 : data_out = 24'b000000001110001010111001;
    16'b0000011111010110 : data_out = 24'b000000001110001011110010;
    16'b0000011111010111 : data_out = 24'b000000001110001100101011;
    16'b0000011111011000 : data_out = 24'b000000001110001101100100;
    16'b0000011111011001 : data_out = 24'b000000001110001110011101;
    16'b0000011111011010 : data_out = 24'b000000001110001111010110;
    16'b0000011111011011 : data_out = 24'b000000001110010000001111;
    16'b0000011111011100 : data_out = 24'b000000001110010001001000;
    16'b0000011111011101 : data_out = 24'b000000001110010010000001;
    16'b0000011111011110 : data_out = 24'b000000001110010010111010;
    16'b0000011111011111 : data_out = 24'b000000001110010011110011;
    16'b0000011111100000 : data_out = 24'b000000001110010100101100;
    16'b0000011111100001 : data_out = 24'b000000001110010101100110;
    16'b0000011111100010 : data_out = 24'b000000001110010110011111;
    16'b0000011111100011 : data_out = 24'b000000001110010111011000;
    16'b0000011111100100 : data_out = 24'b000000001110011000010010;
    16'b0000011111100101 : data_out = 24'b000000001110011001001011;
    16'b0000011111100110 : data_out = 24'b000000001110011010000101;
    16'b0000011111100111 : data_out = 24'b000000001110011010111111;
    16'b0000011111101000 : data_out = 24'b000000001110011011111000;
    16'b0000011111101001 : data_out = 24'b000000001110011100110010;
    16'b0000011111101010 : data_out = 24'b000000001110011101101100;
    16'b0000011111101011 : data_out = 24'b000000001110011110100110;
    16'b0000011111101100 : data_out = 24'b000000001110011111100000;
    16'b0000011111101101 : data_out = 24'b000000001110100000011010;
    16'b0000011111101110 : data_out = 24'b000000001110100001010100;
    16'b0000011111101111 : data_out = 24'b000000001110100010001110;
    16'b0000011111110000 : data_out = 24'b000000001110100011001000;
    16'b0000011111110001 : data_out = 24'b000000001110100100000010;
    16'b0000011111110010 : data_out = 24'b000000001110100100111101;
    16'b0000011111110011 : data_out = 24'b000000001110100101110111;
    16'b0000011111110100 : data_out = 24'b000000001110100110110001;
    16'b0000011111110101 : data_out = 24'b000000001110100111101100;
    16'b0000011111110110 : data_out = 24'b000000001110101000100110;
    16'b0000011111110111 : data_out = 24'b000000001110101001100001;
    16'b0000011111111000 : data_out = 24'b000000001110101010011100;
    16'b0000011111111001 : data_out = 24'b000000001110101011010110;
    16'b0000011111111010 : data_out = 24'b000000001110101100010001;
    16'b0000011111111011 : data_out = 24'b000000001110101101001100;
    16'b0000011111111100 : data_out = 24'b000000001110101110000111;
    16'b0000011111111101 : data_out = 24'b000000001110101111000010;
    16'b0000011111111110 : data_out = 24'b000000001110101111111101;
    16'b0000011111111111 : data_out = 24'b000000001110110000111000;
    16'b0000100000000000 : data_out = 24'b000000001110110001110011;
    16'b0000100000000001 : data_out = 24'b000000001110110010101110;
    16'b0000100000000010 : data_out = 24'b000000001110110011101001;
    16'b0000100000000011 : data_out = 24'b000000001110110100100100;
    16'b0000100000000100 : data_out = 24'b000000001110110101100000;
    16'b0000100000000101 : data_out = 24'b000000001110110110011011;
    16'b0000100000000110 : data_out = 24'b000000001110110111010110;
    16'b0000100000000111 : data_out = 24'b000000001110111000010010;
    16'b0000100000001000 : data_out = 24'b000000001110111001001101;
    16'b0000100000001001 : data_out = 24'b000000001110111010001001;
    16'b0000100000001010 : data_out = 24'b000000001110111011000101;
    16'b0000100000001011 : data_out = 24'b000000001110111100000000;
    16'b0000100000001100 : data_out = 24'b000000001110111100111100;
    16'b0000100000001101 : data_out = 24'b000000001110111101111000;
    16'b0000100000001110 : data_out = 24'b000000001110111110110100;
    16'b0000100000001111 : data_out = 24'b000000001110111111110000;
    16'b0000100000010000 : data_out = 24'b000000001111000000101100;
    16'b0000100000010001 : data_out = 24'b000000001111000001101000;
    16'b0000100000010010 : data_out = 24'b000000001111000010100100;
    16'b0000100000010011 : data_out = 24'b000000001111000011100000;
    16'b0000100000010100 : data_out = 24'b000000001111000100011101;
    16'b0000100000010101 : data_out = 24'b000000001111000101011001;
    16'b0000100000010110 : data_out = 24'b000000001111000110010101;
    16'b0000100000010111 : data_out = 24'b000000001111000111010010;
    16'b0000100000011000 : data_out = 24'b000000001111001000001110;
    16'b0000100000011001 : data_out = 24'b000000001111001001001011;
    16'b0000100000011010 : data_out = 24'b000000001111001010000111;
    16'b0000100000011011 : data_out = 24'b000000001111001011000100;
    16'b0000100000011100 : data_out = 24'b000000001111001100000001;
    16'b0000100000011101 : data_out = 24'b000000001111001100111101;
    16'b0000100000011110 : data_out = 24'b000000001111001101111010;
    16'b0000100000011111 : data_out = 24'b000000001111001110110111;
    16'b0000100000100000 : data_out = 24'b000000001111001111110100;
    16'b0000100000100001 : data_out = 24'b000000001111010000110001;
    16'b0000100000100010 : data_out = 24'b000000001111010001101110;
    16'b0000100000100011 : data_out = 24'b000000001111010010101011;
    16'b0000100000100100 : data_out = 24'b000000001111010011101001;
    16'b0000100000100101 : data_out = 24'b000000001111010100100110;
    16'b0000100000100110 : data_out = 24'b000000001111010101100011;
    16'b0000100000100111 : data_out = 24'b000000001111010110100000;
    16'b0000100000101000 : data_out = 24'b000000001111010111011110;
    16'b0000100000101001 : data_out = 24'b000000001111011000011011;
    16'b0000100000101010 : data_out = 24'b000000001111011001011001;
    16'b0000100000101011 : data_out = 24'b000000001111011010010111;
    16'b0000100000101100 : data_out = 24'b000000001111011011010100;
    16'b0000100000101101 : data_out = 24'b000000001111011100010010;
    16'b0000100000101110 : data_out = 24'b000000001111011101010000;
    16'b0000100000101111 : data_out = 24'b000000001111011110001110;
    16'b0000100000110000 : data_out = 24'b000000001111011111001100;
    16'b0000100000110001 : data_out = 24'b000000001111100000001010;
    16'b0000100000110010 : data_out = 24'b000000001111100001001000;
    16'b0000100000110011 : data_out = 24'b000000001111100010000110;
    16'b0000100000110100 : data_out = 24'b000000001111100011000100;
    16'b0000100000110101 : data_out = 24'b000000001111100100000010;
    16'b0000100000110110 : data_out = 24'b000000001111100101000000;
    16'b0000100000110111 : data_out = 24'b000000001111100101111111;
    16'b0000100000111000 : data_out = 24'b000000001111100110111101;
    16'b0000100000111001 : data_out = 24'b000000001111100111111100;
    16'b0000100000111010 : data_out = 24'b000000001111101000111010;
    16'b0000100000111011 : data_out = 24'b000000001111101001111001;
    16'b0000100000111100 : data_out = 24'b000000001111101010110111;
    16'b0000100000111101 : data_out = 24'b000000001111101011110110;
    16'b0000100000111110 : data_out = 24'b000000001111101100110101;
    16'b0000100000111111 : data_out = 24'b000000001111101101110100;
    16'b0000100001000000 : data_out = 24'b000000001111101110110011;
    16'b0000100001000001 : data_out = 24'b000000001111101111110010;
    16'b0000100001000010 : data_out = 24'b000000001111110000110001;
    16'b0000100001000011 : data_out = 24'b000000001111110001110000;
    16'b0000100001000100 : data_out = 24'b000000001111110010101111;
    16'b0000100001000101 : data_out = 24'b000000001111110011101110;
    16'b0000100001000110 : data_out = 24'b000000001111110100101101;
    16'b0000100001000111 : data_out = 24'b000000001111110101101101;
    16'b0000100001001000 : data_out = 24'b000000001111110110101100;
    16'b0000100001001001 : data_out = 24'b000000001111110111101011;
    16'b0000100001001010 : data_out = 24'b000000001111111000101011;
    16'b0000100001001011 : data_out = 24'b000000001111111001101010;
    16'b0000100001001100 : data_out = 24'b000000001111111010101010;
    16'b0000100001001101 : data_out = 24'b000000001111111011101010;
    16'b0000100001001110 : data_out = 24'b000000001111111100101010;
    16'b0000100001001111 : data_out = 24'b000000001111111101101001;
    16'b0000100001010000 : data_out = 24'b000000001111111110101001;
    16'b0000100001010001 : data_out = 24'b000000001111111111101001;
    16'b0000100001010010 : data_out = 24'b000000010000000000101001;
    16'b0000100001010011 : data_out = 24'b000000010000000001101001;
    16'b0000100001010100 : data_out = 24'b000000010000000010101001;
    16'b0000100001010101 : data_out = 24'b000000010000000011101010;
    16'b0000100001010110 : data_out = 24'b000000010000000100101010;
    16'b0000100001010111 : data_out = 24'b000000010000000101101010;
    16'b0000100001011000 : data_out = 24'b000000010000000110101011;
    16'b0000100001011001 : data_out = 24'b000000010000000111101011;
    16'b0000100001011010 : data_out = 24'b000000010000001000101100;
    16'b0000100001011011 : data_out = 24'b000000010000001001101100;
    16'b0000100001011100 : data_out = 24'b000000010000001010101101;
    16'b0000100001011101 : data_out = 24'b000000010000001011101101;
    16'b0000100001011110 : data_out = 24'b000000010000001100101110;
    16'b0000100001011111 : data_out = 24'b000000010000001101101111;
    16'b0000100001100000 : data_out = 24'b000000010000001110110000;
    16'b0000100001100001 : data_out = 24'b000000010000001111110001;
    16'b0000100001100010 : data_out = 24'b000000010000010000110010;
    16'b0000100001100011 : data_out = 24'b000000010000010001110011;
    16'b0000100001100100 : data_out = 24'b000000010000010010110100;
    16'b0000100001100101 : data_out = 24'b000000010000010011110101;
    16'b0000100001100110 : data_out = 24'b000000010000010100110111;
    16'b0000100001100111 : data_out = 24'b000000010000010101111000;
    16'b0000100001101000 : data_out = 24'b000000010000010110111001;
    16'b0000100001101001 : data_out = 24'b000000010000010111111011;
    16'b0000100001101010 : data_out = 24'b000000010000011000111100;
    16'b0000100001101011 : data_out = 24'b000000010000011001111110;
    16'b0000100001101100 : data_out = 24'b000000010000011011000000;
    16'b0000100001101101 : data_out = 24'b000000010000011100000001;
    16'b0000100001101110 : data_out = 24'b000000010000011101000011;
    16'b0000100001101111 : data_out = 24'b000000010000011110000101;
    16'b0000100001110000 : data_out = 24'b000000010000011111000111;
    16'b0000100001110001 : data_out = 24'b000000010000100000001001;
    16'b0000100001110010 : data_out = 24'b000000010000100001001011;
    16'b0000100001110011 : data_out = 24'b000000010000100010001101;
    16'b0000100001110100 : data_out = 24'b000000010000100011001111;
    16'b0000100001110101 : data_out = 24'b000000010000100100010001;
    16'b0000100001110110 : data_out = 24'b000000010000100101010100;
    16'b0000100001110111 : data_out = 24'b000000010000100110010110;
    16'b0000100001111000 : data_out = 24'b000000010000100111011000;
    16'b0000100001111001 : data_out = 24'b000000010000101000011011;
    16'b0000100001111010 : data_out = 24'b000000010000101001011110;
    16'b0000100001111011 : data_out = 24'b000000010000101010100000;
    16'b0000100001111100 : data_out = 24'b000000010000101011100011;
    16'b0000100001111101 : data_out = 24'b000000010000101100100110;
    16'b0000100001111110 : data_out = 24'b000000010000101101101000;
    16'b0000100001111111 : data_out = 24'b000000010000101110101011;
    16'b0000100010000000 : data_out = 24'b000000010000101111101110;
    16'b0000100010000001 : data_out = 24'b000000010000110000110001;
    16'b0000100010000010 : data_out = 24'b000000010000110001110100;
    16'b0000100010000011 : data_out = 24'b000000010000110010111000;
    16'b0000100010000100 : data_out = 24'b000000010000110011111011;
    16'b0000100010000101 : data_out = 24'b000000010000110100111110;
    16'b0000100010000110 : data_out = 24'b000000010000110110000001;
    16'b0000100010000111 : data_out = 24'b000000010000110111000101;
    16'b0000100010001000 : data_out = 24'b000000010000111000001000;
    16'b0000100010001001 : data_out = 24'b000000010000111001001100;
    16'b0000100010001010 : data_out = 24'b000000010000111010001111;
    16'b0000100010001011 : data_out = 24'b000000010000111011010011;
    16'b0000100010001100 : data_out = 24'b000000010000111100010111;
    16'b0000100010001101 : data_out = 24'b000000010000111101011011;
    16'b0000100010001110 : data_out = 24'b000000010000111110011110;
    16'b0000100010001111 : data_out = 24'b000000010000111111100010;
    16'b0000100010010000 : data_out = 24'b000000010001000000100110;
    16'b0000100010010001 : data_out = 24'b000000010001000001101010;
    16'b0000100010010010 : data_out = 24'b000000010001000010101111;
    16'b0000100010010011 : data_out = 24'b000000010001000011110011;
    16'b0000100010010100 : data_out = 24'b000000010001000100110111;
    16'b0000100010010101 : data_out = 24'b000000010001000101111011;
    16'b0000100010010110 : data_out = 24'b000000010001000111000000;
    16'b0000100010010111 : data_out = 24'b000000010001001000000100;
    16'b0000100010011000 : data_out = 24'b000000010001001001001001;
    16'b0000100010011001 : data_out = 24'b000000010001001010001101;
    16'b0000100010011010 : data_out = 24'b000000010001001011010010;
    16'b0000100010011011 : data_out = 24'b000000010001001100010111;
    16'b0000100010011100 : data_out = 24'b000000010001001101011100;
    16'b0000100010011101 : data_out = 24'b000000010001001110100001;
    16'b0000100010011110 : data_out = 24'b000000010001001111100101;
    16'b0000100010011111 : data_out = 24'b000000010001010000101011;
    16'b0000100010100000 : data_out = 24'b000000010001010001110000;
    16'b0000100010100001 : data_out = 24'b000000010001010010110101;
    16'b0000100010100010 : data_out = 24'b000000010001010011111010;
    16'b0000100010100011 : data_out = 24'b000000010001010100111111;
    16'b0000100010100100 : data_out = 24'b000000010001010110000101;
    16'b0000100010100101 : data_out = 24'b000000010001010111001010;
    16'b0000100010100110 : data_out = 24'b000000010001011000001111;
    16'b0000100010100111 : data_out = 24'b000000010001011001010101;
    16'b0000100010101000 : data_out = 24'b000000010001011010011011;
    16'b0000100010101001 : data_out = 24'b000000010001011011100000;
    16'b0000100010101010 : data_out = 24'b000000010001011100100110;
    16'b0000100010101011 : data_out = 24'b000000010001011101101100;
    16'b0000100010101100 : data_out = 24'b000000010001011110110010;
    16'b0000100010101101 : data_out = 24'b000000010001011111111000;
    16'b0000100010101110 : data_out = 24'b000000010001100000111110;
    16'b0000100010101111 : data_out = 24'b000000010001100010000100;
    16'b0000100010110000 : data_out = 24'b000000010001100011001010;
    16'b0000100010110001 : data_out = 24'b000000010001100100010000;
    16'b0000100010110010 : data_out = 24'b000000010001100101010111;
    16'b0000100010110011 : data_out = 24'b000000010001100110011101;
    16'b0000100010110100 : data_out = 24'b000000010001100111100011;
    16'b0000100010110101 : data_out = 24'b000000010001101000101010;
    16'b0000100010110110 : data_out = 24'b000000010001101001110000;
    16'b0000100010110111 : data_out = 24'b000000010001101010110111;
    16'b0000100010111000 : data_out = 24'b000000010001101011111110;
    16'b0000100010111001 : data_out = 24'b000000010001101101000101;
    16'b0000100010111010 : data_out = 24'b000000010001101110001011;
    16'b0000100010111011 : data_out = 24'b000000010001101111010010;
    16'b0000100010111100 : data_out = 24'b000000010001110000011001;
    16'b0000100010111101 : data_out = 24'b000000010001110001100000;
    16'b0000100010111110 : data_out = 24'b000000010001110010101000;
    16'b0000100010111111 : data_out = 24'b000000010001110011101111;
    16'b0000100011000000 : data_out = 24'b000000010001110100110110;
    16'b0000100011000001 : data_out = 24'b000000010001110101111101;
    16'b0000100011000010 : data_out = 24'b000000010001110111000101;
    16'b0000100011000011 : data_out = 24'b000000010001111000001100;
    16'b0000100011000100 : data_out = 24'b000000010001111001010100;
    16'b0000100011000101 : data_out = 24'b000000010001111010011011;
    16'b0000100011000110 : data_out = 24'b000000010001111011100011;
    16'b0000100011000111 : data_out = 24'b000000010001111100101011;
    16'b0000100011001000 : data_out = 24'b000000010001111101110011;
    16'b0000100011001001 : data_out = 24'b000000010001111110111011;
    16'b0000100011001010 : data_out = 24'b000000010010000000000011;
    16'b0000100011001011 : data_out = 24'b000000010010000001001011;
    16'b0000100011001100 : data_out = 24'b000000010010000010010011;
    16'b0000100011001101 : data_out = 24'b000000010010000011011011;
    16'b0000100011001110 : data_out = 24'b000000010010000100100011;
    16'b0000100011001111 : data_out = 24'b000000010010000101101011;
    16'b0000100011010000 : data_out = 24'b000000010010000110110100;
    16'b0000100011010001 : data_out = 24'b000000010010000111111100;
    16'b0000100011010010 : data_out = 24'b000000010010001001000101;
    16'b0000100011010011 : data_out = 24'b000000010010001010001101;
    16'b0000100011010100 : data_out = 24'b000000010010001011010110;
    16'b0000100011010101 : data_out = 24'b000000010010001100011111;
    16'b0000100011010110 : data_out = 24'b000000010010001101101000;
    16'b0000100011010111 : data_out = 24'b000000010010001110110001;
    16'b0000100011011000 : data_out = 24'b000000010010001111111001;
    16'b0000100011011001 : data_out = 24'b000000010010010001000011;
    16'b0000100011011010 : data_out = 24'b000000010010010010001100;
    16'b0000100011011011 : data_out = 24'b000000010010010011010101;
    16'b0000100011011100 : data_out = 24'b000000010010010100011110;
    16'b0000100011011101 : data_out = 24'b000000010010010101100111;
    16'b0000100011011110 : data_out = 24'b000000010010010110110001;
    16'b0000100011011111 : data_out = 24'b000000010010010111111010;
    16'b0000100011100000 : data_out = 24'b000000010010011001000100;
    16'b0000100011100001 : data_out = 24'b000000010010011010001101;
    16'b0000100011100010 : data_out = 24'b000000010010011011010111;
    16'b0000100011100011 : data_out = 24'b000000010010011100100001;
    16'b0000100011100100 : data_out = 24'b000000010010011101101011;
    16'b0000100011100101 : data_out = 24'b000000010010011110110100;
    16'b0000100011100110 : data_out = 24'b000000010010011111111110;
    16'b0000100011100111 : data_out = 24'b000000010010100001001000;
    16'b0000100011101000 : data_out = 24'b000000010010100010010011;
    16'b0000100011101001 : data_out = 24'b000000010010100011011101;
    16'b0000100011101010 : data_out = 24'b000000010010100100100111;
    16'b0000100011101011 : data_out = 24'b000000010010100101110001;
    16'b0000100011101100 : data_out = 24'b000000010010100110111100;
    16'b0000100011101101 : data_out = 24'b000000010010101000000110;
    16'b0000100011101110 : data_out = 24'b000000010010101001010001;
    16'b0000100011101111 : data_out = 24'b000000010010101010011011;
    16'b0000100011110000 : data_out = 24'b000000010010101011100110;
    16'b0000100011110001 : data_out = 24'b000000010010101100110001;
    16'b0000100011110010 : data_out = 24'b000000010010101101111100;
    16'b0000100011110011 : data_out = 24'b000000010010101111000111;
    16'b0000100011110100 : data_out = 24'b000000010010110000010010;
    16'b0000100011110101 : data_out = 24'b000000010010110001011101;
    16'b0000100011110110 : data_out = 24'b000000010010110010101000;
    16'b0000100011110111 : data_out = 24'b000000010010110011110011;
    16'b0000100011111000 : data_out = 24'b000000010010110100111110;
    16'b0000100011111001 : data_out = 24'b000000010010110110001010;
    16'b0000100011111010 : data_out = 24'b000000010010110111010101;
    16'b0000100011111011 : data_out = 24'b000000010010111000100000;
    16'b0000100011111100 : data_out = 24'b000000010010111001101100;
    16'b0000100011111101 : data_out = 24'b000000010010111010111000;
    16'b0000100011111110 : data_out = 24'b000000010010111100000011;
    16'b0000100011111111 : data_out = 24'b000000010010111101001111;
    16'b0000100100000000 : data_out = 24'b000000010010111110011011;
    16'b0000100100000001 : data_out = 24'b000000010010111111100111;
    16'b0000100100000010 : data_out = 24'b000000010011000000110011;
    16'b0000100100000011 : data_out = 24'b000000010011000001111111;
    16'b0000100100000100 : data_out = 24'b000000010011000011001011;
    16'b0000100100000101 : data_out = 24'b000000010011000100010111;
    16'b0000100100000110 : data_out = 24'b000000010011000101100100;
    16'b0000100100000111 : data_out = 24'b000000010011000110110000;
    16'b0000100100001000 : data_out = 24'b000000010011000111111101;
    16'b0000100100001001 : data_out = 24'b000000010011001001001001;
    16'b0000100100001010 : data_out = 24'b000000010011001010010110;
    16'b0000100100001011 : data_out = 24'b000000010011001011100010;
    16'b0000100100001100 : data_out = 24'b000000010011001100101111;
    16'b0000100100001101 : data_out = 24'b000000010011001101111100;
    16'b0000100100001110 : data_out = 24'b000000010011001111001001;
    16'b0000100100001111 : data_out = 24'b000000010011010000010110;
    16'b0000100100010000 : data_out = 24'b000000010011010001100011;
    16'b0000100100010001 : data_out = 24'b000000010011010010110000;
    16'b0000100100010010 : data_out = 24'b000000010011010011111101;
    16'b0000100100010011 : data_out = 24'b000000010011010101001011;
    16'b0000100100010100 : data_out = 24'b000000010011010110011000;
    16'b0000100100010101 : data_out = 24'b000000010011010111100101;
    16'b0000100100010110 : data_out = 24'b000000010011011000110011;
    16'b0000100100010111 : data_out = 24'b000000010011011010000001;
    16'b0000100100011000 : data_out = 24'b000000010011011011001110;
    16'b0000100100011001 : data_out = 24'b000000010011011100011100;
    16'b0000100100011010 : data_out = 24'b000000010011011101101010;
    16'b0000100100011011 : data_out = 24'b000000010011011110111000;
    16'b0000100100011100 : data_out = 24'b000000010011100000000110;
    16'b0000100100011101 : data_out = 24'b000000010011100001010100;
    16'b0000100100011110 : data_out = 24'b000000010011100010100010;
    16'b0000100100011111 : data_out = 24'b000000010011100011110000;
    16'b0000100100100000 : data_out = 24'b000000010011100100111110;
    16'b0000100100100001 : data_out = 24'b000000010011100110001101;
    16'b0000100100100010 : data_out = 24'b000000010011100111011011;
    16'b0000100100100011 : data_out = 24'b000000010011101000101010;
    16'b0000100100100100 : data_out = 24'b000000010011101001111000;
    16'b0000100100100101 : data_out = 24'b000000010011101011000111;
    16'b0000100100100110 : data_out = 24'b000000010011101100010101;
    16'b0000100100100111 : data_out = 24'b000000010011101101100100;
    16'b0000100100101000 : data_out = 24'b000000010011101110110011;
    16'b0000100100101001 : data_out = 24'b000000010011110000000010;
    16'b0000100100101010 : data_out = 24'b000000010011110001010001;
    16'b0000100100101011 : data_out = 24'b000000010011110010100000;
    16'b0000100100101100 : data_out = 24'b000000010011110011110000;
    16'b0000100100101101 : data_out = 24'b000000010011110100111111;
    16'b0000100100101110 : data_out = 24'b000000010011110110001110;
    16'b0000100100101111 : data_out = 24'b000000010011110111011110;
    16'b0000100100110000 : data_out = 24'b000000010011111000101101;
    16'b0000100100110001 : data_out = 24'b000000010011111001111101;
    16'b0000100100110010 : data_out = 24'b000000010011111011001100;
    16'b0000100100110011 : data_out = 24'b000000010011111100011100;
    16'b0000100100110100 : data_out = 24'b000000010011111101101100;
    16'b0000100100110101 : data_out = 24'b000000010011111110111100;
    16'b0000100100110110 : data_out = 24'b000000010100000000001100;
    16'b0000100100110111 : data_out = 24'b000000010100000001011100;
    16'b0000100100111000 : data_out = 24'b000000010100000010101100;
    16'b0000100100111001 : data_out = 24'b000000010100000011111100;
    16'b0000100100111010 : data_out = 24'b000000010100000101001100;
    16'b0000100100111011 : data_out = 24'b000000010100000110011101;
    16'b0000100100111100 : data_out = 24'b000000010100000111101101;
    16'b0000100100111101 : data_out = 24'b000000010100001000111110;
    16'b0000100100111110 : data_out = 24'b000000010100001010001110;
    16'b0000100100111111 : data_out = 24'b000000010100001011011111;
    16'b0000100101000000 : data_out = 24'b000000010100001100110000;
    16'b0000100101000001 : data_out = 24'b000000010100001110000001;
    16'b0000100101000010 : data_out = 24'b000000010100001111010010;
    16'b0000100101000011 : data_out = 24'b000000010100010000100011;
    16'b0000100101000100 : data_out = 24'b000000010100010001110100;
    16'b0000100101000101 : data_out = 24'b000000010100010011000101;
    16'b0000100101000110 : data_out = 24'b000000010100010100010110;
    16'b0000100101000111 : data_out = 24'b000000010100010101100111;
    16'b0000100101001000 : data_out = 24'b000000010100010110111001;
    16'b0000100101001001 : data_out = 24'b000000010100011000001010;
    16'b0000100101001010 : data_out = 24'b000000010100011001011100;
    16'b0000100101001011 : data_out = 24'b000000010100011010101101;
    16'b0000100101001100 : data_out = 24'b000000010100011011111111;
    16'b0000100101001101 : data_out = 24'b000000010100011101010001;
    16'b0000100101001110 : data_out = 24'b000000010100011110100011;
    16'b0000100101001111 : data_out = 24'b000000010100011111110101;
    16'b0000100101010000 : data_out = 24'b000000010100100001000111;
    16'b0000100101010001 : data_out = 24'b000000010100100010011001;
    16'b0000100101010010 : data_out = 24'b000000010100100011101011;
    16'b0000100101010011 : data_out = 24'b000000010100100100111101;
    16'b0000100101010100 : data_out = 24'b000000010100100110010000;
    16'b0000100101010101 : data_out = 24'b000000010100100111100010;
    16'b0000100101010110 : data_out = 24'b000000010100101000110101;
    16'b0000100101010111 : data_out = 24'b000000010100101010000111;
    16'b0000100101011000 : data_out = 24'b000000010100101011011010;
    16'b0000100101011001 : data_out = 24'b000000010100101100101101;
    16'b0000100101011010 : data_out = 24'b000000010100101101111111;
    16'b0000100101011011 : data_out = 24'b000000010100101111010010;
    16'b0000100101011100 : data_out = 24'b000000010100110000100101;
    16'b0000100101011101 : data_out = 24'b000000010100110001111000;
    16'b0000100101011110 : data_out = 24'b000000010100110011001100;
    16'b0000100101011111 : data_out = 24'b000000010100110100011111;
    16'b0000100101100000 : data_out = 24'b000000010100110101110010;
    16'b0000100101100001 : data_out = 24'b000000010100110111000110;
    16'b0000100101100010 : data_out = 24'b000000010100111000011001;
    16'b0000100101100011 : data_out = 24'b000000010100111001101101;
    16'b0000100101100100 : data_out = 24'b000000010100111011000000;
    16'b0000100101100101 : data_out = 24'b000000010100111100010100;
    16'b0000100101100110 : data_out = 24'b000000010100111101101000;
    16'b0000100101100111 : data_out = 24'b000000010100111110111100;
    16'b0000100101101000 : data_out = 24'b000000010101000000010000;
    16'b0000100101101001 : data_out = 24'b000000010101000001100100;
    16'b0000100101101010 : data_out = 24'b000000010101000010111000;
    16'b0000100101101011 : data_out = 24'b000000010101000100001100;
    16'b0000100101101100 : data_out = 24'b000000010101000101100000;
    16'b0000100101101101 : data_out = 24'b000000010101000110110101;
    16'b0000100101101110 : data_out = 24'b000000010101001000001001;
    16'b0000100101101111 : data_out = 24'b000000010101001001011110;
    16'b0000100101110000 : data_out = 24'b000000010101001010110010;
    16'b0000100101110001 : data_out = 24'b000000010101001100000111;
    16'b0000100101110010 : data_out = 24'b000000010101001101011100;
    16'b0000100101110011 : data_out = 24'b000000010101001110110001;
    16'b0000100101110100 : data_out = 24'b000000010101010000000110;
    16'b0000100101110101 : data_out = 24'b000000010101010001011011;
    16'b0000100101110110 : data_out = 24'b000000010101010010110000;
    16'b0000100101110111 : data_out = 24'b000000010101010100000101;
    16'b0000100101111000 : data_out = 24'b000000010101010101011010;
    16'b0000100101111001 : data_out = 24'b000000010101010110110000;
    16'b0000100101111010 : data_out = 24'b000000010101011000000101;
    16'b0000100101111011 : data_out = 24'b000000010101011001011011;
    16'b0000100101111100 : data_out = 24'b000000010101011010110000;
    16'b0000100101111101 : data_out = 24'b000000010101011100000110;
    16'b0000100101111110 : data_out = 24'b000000010101011101011100;
    16'b0000100101111111 : data_out = 24'b000000010101011110110010;
    16'b0000100110000000 : data_out = 24'b000000010101100000001000;
    16'b0000100110000001 : data_out = 24'b000000010101100001011110;
    16'b0000100110000010 : data_out = 24'b000000010101100010110100;
    16'b0000100110000011 : data_out = 24'b000000010101100100001010;
    16'b0000100110000100 : data_out = 24'b000000010101100101100001;
    16'b0000100110000101 : data_out = 24'b000000010101100110110111;
    16'b0000100110000110 : data_out = 24'b000000010101101000001101;
    16'b0000100110000111 : data_out = 24'b000000010101101001100100;
    16'b0000100110001000 : data_out = 24'b000000010101101010111011;
    16'b0000100110001001 : data_out = 24'b000000010101101100010001;
    16'b0000100110001010 : data_out = 24'b000000010101101101101000;
    16'b0000100110001011 : data_out = 24'b000000010101101110111111;
    16'b0000100110001100 : data_out = 24'b000000010101110000010110;
    16'b0000100110001101 : data_out = 24'b000000010101110001101101;
    16'b0000100110001110 : data_out = 24'b000000010101110011000100;
    16'b0000100110001111 : data_out = 24'b000000010101110100011011;
    16'b0000100110010000 : data_out = 24'b000000010101110101110011;
    16'b0000100110010001 : data_out = 24'b000000010101110111001010;
    16'b0000100110010010 : data_out = 24'b000000010101111000100010;
    16'b0000100110010011 : data_out = 24'b000000010101111001111001;
    16'b0000100110010100 : data_out = 24'b000000010101111011010001;
    16'b0000100110010101 : data_out = 24'b000000010101111100101001;
    16'b0000100110010110 : data_out = 24'b000000010101111110000000;
    16'b0000100110010111 : data_out = 24'b000000010101111111011000;
    16'b0000100110011000 : data_out = 24'b000000010110000000110000;
    16'b0000100110011001 : data_out = 24'b000000010110000010001000;
    16'b0000100110011010 : data_out = 24'b000000010110000011100001;
    16'b0000100110011011 : data_out = 24'b000000010110000100111001;
    16'b0000100110011100 : data_out = 24'b000000010110000110010001;
    16'b0000100110011101 : data_out = 24'b000000010110000111101010;
    16'b0000100110011110 : data_out = 24'b000000010110001001000010;
    16'b0000100110011111 : data_out = 24'b000000010110001010011011;
    16'b0000100110100000 : data_out = 24'b000000010110001011110100;
    16'b0000100110100001 : data_out = 24'b000000010110001101001100;
    16'b0000100110100010 : data_out = 24'b000000010110001110100101;
    16'b0000100110100011 : data_out = 24'b000000010110001111111110;
    16'b0000100110100100 : data_out = 24'b000000010110010001010111;
    16'b0000100110100101 : data_out = 24'b000000010110010010110000;
    16'b0000100110100110 : data_out = 24'b000000010110010100001010;
    16'b0000100110100111 : data_out = 24'b000000010110010101100011;
    16'b0000100110101000 : data_out = 24'b000000010110010110111100;
    16'b0000100110101001 : data_out = 24'b000000010110011000010110;
    16'b0000100110101010 : data_out = 24'b000000010110011001101111;
    16'b0000100110101011 : data_out = 24'b000000010110011011001001;
    16'b0000100110101100 : data_out = 24'b000000010110011100100011;
    16'b0000100110101101 : data_out = 24'b000000010110011101111100;
    16'b0000100110101110 : data_out = 24'b000000010110011111010110;
    16'b0000100110101111 : data_out = 24'b000000010110100000110000;
    16'b0000100110110000 : data_out = 24'b000000010110100010001010;
    16'b0000100110110001 : data_out = 24'b000000010110100011100101;
    16'b0000100110110010 : data_out = 24'b000000010110100100111111;
    16'b0000100110110011 : data_out = 24'b000000010110100110011001;
    16'b0000100110110100 : data_out = 24'b000000010110100111110100;
    16'b0000100110110101 : data_out = 24'b000000010110101001001110;
    16'b0000100110110110 : data_out = 24'b000000010110101010101001;
    16'b0000100110110111 : data_out = 24'b000000010110101100000100;
    16'b0000100110111000 : data_out = 24'b000000010110101101011110;
    16'b0000100110111001 : data_out = 24'b000000010110101110111001;
    16'b0000100110111010 : data_out = 24'b000000010110110000010100;
    16'b0000100110111011 : data_out = 24'b000000010110110001101111;
    16'b0000100110111100 : data_out = 24'b000000010110110011001010;
    16'b0000100110111101 : data_out = 24'b000000010110110100100110;
    16'b0000100110111110 : data_out = 24'b000000010110110110000001;
    16'b0000100110111111 : data_out = 24'b000000010110110111011100;
    16'b0000100111000000 : data_out = 24'b000000010110111000111000;
    16'b0000100111000001 : data_out = 24'b000000010110111010010100;
    16'b0000100111000010 : data_out = 24'b000000010110111011101111;
    16'b0000100111000011 : data_out = 24'b000000010110111101001011;
    16'b0000100111000100 : data_out = 24'b000000010110111110100111;
    16'b0000100111000101 : data_out = 24'b000000010111000000000011;
    16'b0000100111000110 : data_out = 24'b000000010111000001011111;
    16'b0000100111000111 : data_out = 24'b000000010111000010111011;
    16'b0000100111001000 : data_out = 24'b000000010111000100010111;
    16'b0000100111001001 : data_out = 24'b000000010111000101110100;
    16'b0000100111001010 : data_out = 24'b000000010111000111010000;
    16'b0000100111001011 : data_out = 24'b000000010111001000101101;
    16'b0000100111001100 : data_out = 24'b000000010111001010001001;
    16'b0000100111001101 : data_out = 24'b000000010111001011100110;
    16'b0000100111001110 : data_out = 24'b000000010111001101000011;
    16'b0000100111001111 : data_out = 24'b000000010111001110011111;
    16'b0000100111010000 : data_out = 24'b000000010111001111111100;
    16'b0000100111010001 : data_out = 24'b000000010111010001011001;
    16'b0000100111010010 : data_out = 24'b000000010111010010110111;
    16'b0000100111010011 : data_out = 24'b000000010111010100010100;
    16'b0000100111010100 : data_out = 24'b000000010111010101110001;
    16'b0000100111010101 : data_out = 24'b000000010111010111001110;
    16'b0000100111010110 : data_out = 24'b000000010111011000101100;
    16'b0000100111010111 : data_out = 24'b000000010111011010001010;
    16'b0000100111011000 : data_out = 24'b000000010111011011100111;
    16'b0000100111011001 : data_out = 24'b000000010111011101000101;
    16'b0000100111011010 : data_out = 24'b000000010111011110100011;
    16'b0000100111011011 : data_out = 24'b000000010111100000000001;
    16'b0000100111011100 : data_out = 24'b000000010111100001011111;
    16'b0000100111011101 : data_out = 24'b000000010111100010111101;
    16'b0000100111011110 : data_out = 24'b000000010111100100011011;
    16'b0000100111011111 : data_out = 24'b000000010111100101111010;
    16'b0000100111100000 : data_out = 24'b000000010111100111011000;
    16'b0000100111100001 : data_out = 24'b000000010111101000110111;
    16'b0000100111100010 : data_out = 24'b000000010111101010010101;
    16'b0000100111100011 : data_out = 24'b000000010111101011110100;
    16'b0000100111100100 : data_out = 24'b000000010111101101010011;
    16'b0000100111100101 : data_out = 24'b000000010111101110110001;
    16'b0000100111100110 : data_out = 24'b000000010111110000010000;
    16'b0000100111100111 : data_out = 24'b000000010111110001101111;
    16'b0000100111101000 : data_out = 24'b000000010111110011001111;
    16'b0000100111101001 : data_out = 24'b000000010111110100101110;
    16'b0000100111101010 : data_out = 24'b000000010111110110001101;
    16'b0000100111101011 : data_out = 24'b000000010111110111101101;
    16'b0000100111101100 : data_out = 24'b000000010111111001001100;
    16'b0000100111101101 : data_out = 24'b000000010111111010101100;
    16'b0000100111101110 : data_out = 24'b000000010111111100001100;
    16'b0000100111101111 : data_out = 24'b000000010111111101101011;
    16'b0000100111110000 : data_out = 24'b000000010111111111001011;
    16'b0000100111110001 : data_out = 24'b000000011000000000101011;
    16'b0000100111110010 : data_out = 24'b000000011000000010001011;
    16'b0000100111110011 : data_out = 24'b000000011000000011101100;
    16'b0000100111110100 : data_out = 24'b000000011000000101001100;
    16'b0000100111110101 : data_out = 24'b000000011000000110101100;
    16'b0000100111110110 : data_out = 24'b000000011000001000001101;
    16'b0000100111110111 : data_out = 24'b000000011000001001101101;
    16'b0000100111111000 : data_out = 24'b000000011000001011001110;
    16'b0000100111111001 : data_out = 24'b000000011000001100101111;
    16'b0000100111111010 : data_out = 24'b000000011000001110001111;
    16'b0000100111111011 : data_out = 24'b000000011000001111110000;
    16'b0000100111111100 : data_out = 24'b000000011000010001010001;
    16'b0000100111111101 : data_out = 24'b000000011000010010110011;
    16'b0000100111111110 : data_out = 24'b000000011000010100010100;
    16'b0000100111111111 : data_out = 24'b000000011000010101110101;
    16'b0000101000000000 : data_out = 24'b000000011000010111010110;
    16'b0000101000000001 : data_out = 24'b000000011000011000111000;
    16'b0000101000000010 : data_out = 24'b000000011000011010011010;
    16'b0000101000000011 : data_out = 24'b000000011000011011111011;
    16'b0000101000000100 : data_out = 24'b000000011000011101011101;
    16'b0000101000000101 : data_out = 24'b000000011000011110111111;
    16'b0000101000000110 : data_out = 24'b000000011000100000100001;
    16'b0000101000000111 : data_out = 24'b000000011000100010000011;
    16'b0000101000001000 : data_out = 24'b000000011000100011100101;
    16'b0000101000001001 : data_out = 24'b000000011000100101000111;
    16'b0000101000001010 : data_out = 24'b000000011000100110101010;
    16'b0000101000001011 : data_out = 24'b000000011000101000001100;
    16'b0000101000001100 : data_out = 24'b000000011000101001101111;
    16'b0000101000001101 : data_out = 24'b000000011000101011010010;
    16'b0000101000001110 : data_out = 24'b000000011000101100110100;
    16'b0000101000001111 : data_out = 24'b000000011000101110010111;
    16'b0000101000010000 : data_out = 24'b000000011000101111111010;
    16'b0000101000010001 : data_out = 24'b000000011000110001011101;
    16'b0000101000010010 : data_out = 24'b000000011000110011000000;
    16'b0000101000010011 : data_out = 24'b000000011000110100100100;
    16'b0000101000010100 : data_out = 24'b000000011000110110000111;
    16'b0000101000010101 : data_out = 24'b000000011000110111101010;
    16'b0000101000010110 : data_out = 24'b000000011000111001001110;
    16'b0000101000010111 : data_out = 24'b000000011000111010110001;
    16'b0000101000011000 : data_out = 24'b000000011000111100010101;
    16'b0000101000011001 : data_out = 24'b000000011000111101111001;
    16'b0000101000011010 : data_out = 24'b000000011000111111011101;
    16'b0000101000011011 : data_out = 24'b000000011001000001000001;
    16'b0000101000011100 : data_out = 24'b000000011001000010100101;
    16'b0000101000011101 : data_out = 24'b000000011001000100001001;
    16'b0000101000011110 : data_out = 24'b000000011001000101101110;
    16'b0000101000011111 : data_out = 24'b000000011001000111010010;
    16'b0000101000100000 : data_out = 24'b000000011001001000110110;
    16'b0000101000100001 : data_out = 24'b000000011001001010011011;
    16'b0000101000100010 : data_out = 24'b000000011001001100000000;
    16'b0000101000100011 : data_out = 24'b000000011001001101100101;
    16'b0000101000100100 : data_out = 24'b000000011001001111001001;
    16'b0000101000100101 : data_out = 24'b000000011001010000101110;
    16'b0000101000100110 : data_out = 24'b000000011001010010010100;
    16'b0000101000100111 : data_out = 24'b000000011001010011111001;
    16'b0000101000101000 : data_out = 24'b000000011001010101011110;
    16'b0000101000101001 : data_out = 24'b000000011001010111000011;
    16'b0000101000101010 : data_out = 24'b000000011001011000101001;
    16'b0000101000101011 : data_out = 24'b000000011001011010001111;
    16'b0000101000101100 : data_out = 24'b000000011001011011110100;
    16'b0000101000101101 : data_out = 24'b000000011001011101011010;
    16'b0000101000101110 : data_out = 24'b000000011001011111000000;
    16'b0000101000101111 : data_out = 24'b000000011001100000100110;
    16'b0000101000110000 : data_out = 24'b000000011001100010001100;
    16'b0000101000110001 : data_out = 24'b000000011001100011110010;
    16'b0000101000110010 : data_out = 24'b000000011001100101011000;
    16'b0000101000110011 : data_out = 24'b000000011001100110111111;
    16'b0000101000110100 : data_out = 24'b000000011001101000100101;
    16'b0000101000110101 : data_out = 24'b000000011001101010001100;
    16'b0000101000110110 : data_out = 24'b000000011001101011110011;
    16'b0000101000110111 : data_out = 24'b000000011001101101011001;
    16'b0000101000111000 : data_out = 24'b000000011001101111000000;
    16'b0000101000111001 : data_out = 24'b000000011001110000100111;
    16'b0000101000111010 : data_out = 24'b000000011001110010001110;
    16'b0000101000111011 : data_out = 24'b000000011001110011110110;
    16'b0000101000111100 : data_out = 24'b000000011001110101011101;
    16'b0000101000111101 : data_out = 24'b000000011001110111000100;
    16'b0000101000111110 : data_out = 24'b000000011001111000101100;
    16'b0000101000111111 : data_out = 24'b000000011001111010010011;
    16'b0000101001000000 : data_out = 24'b000000011001111011111011;
    16'b0000101001000001 : data_out = 24'b000000011001111101100011;
    16'b0000101001000010 : data_out = 24'b000000011001111111001011;
    16'b0000101001000011 : data_out = 24'b000000011010000000110011;
    16'b0000101001000100 : data_out = 24'b000000011010000010011011;
    16'b0000101001000101 : data_out = 24'b000000011010000100000011;
    16'b0000101001000110 : data_out = 24'b000000011010000101101011;
    16'b0000101001000111 : data_out = 24'b000000011010000111010100;
    16'b0000101001001000 : data_out = 24'b000000011010001000111100;
    16'b0000101001001001 : data_out = 24'b000000011010001010100101;
    16'b0000101001001010 : data_out = 24'b000000011010001100001110;
    16'b0000101001001011 : data_out = 24'b000000011010001101110110;
    16'b0000101001001100 : data_out = 24'b000000011010001111011111;
    16'b0000101001001101 : data_out = 24'b000000011010010001001000;
    16'b0000101001001110 : data_out = 24'b000000011010010010110001;
    16'b0000101001001111 : data_out = 24'b000000011010010100011011;
    16'b0000101001010000 : data_out = 24'b000000011010010110000100;
    16'b0000101001010001 : data_out = 24'b000000011010010111101101;
    16'b0000101001010010 : data_out = 24'b000000011010011001010111;
    16'b0000101001010011 : data_out = 24'b000000011010011011000001;
    16'b0000101001010100 : data_out = 24'b000000011010011100101010;
    16'b0000101001010101 : data_out = 24'b000000011010011110010100;
    16'b0000101001010110 : data_out = 24'b000000011010011111111110;
    16'b0000101001010111 : data_out = 24'b000000011010100001101000;
    16'b0000101001011000 : data_out = 24'b000000011010100011010010;
    16'b0000101001011001 : data_out = 24'b000000011010100100111101;
    16'b0000101001011010 : data_out = 24'b000000011010100110100111;
    16'b0000101001011011 : data_out = 24'b000000011010101000010001;
    16'b0000101001011100 : data_out = 24'b000000011010101001111100;
    16'b0000101001011101 : data_out = 24'b000000011010101011100111;
    16'b0000101001011110 : data_out = 24'b000000011010101101010001;
    16'b0000101001011111 : data_out = 24'b000000011010101110111100;
    16'b0000101001100000 : data_out = 24'b000000011010110000100111;
    16'b0000101001100001 : data_out = 24'b000000011010110010010010;
    16'b0000101001100010 : data_out = 24'b000000011010110011111110;
    16'b0000101001100011 : data_out = 24'b000000011010110101101001;
    16'b0000101001100100 : data_out = 24'b000000011010110111010100;
    16'b0000101001100101 : data_out = 24'b000000011010111001000000;
    16'b0000101001100110 : data_out = 24'b000000011010111010101011;
    16'b0000101001100111 : data_out = 24'b000000011010111100010111;
    16'b0000101001101000 : data_out = 24'b000000011010111110000011;
    16'b0000101001101001 : data_out = 24'b000000011010111111101111;
    16'b0000101001101010 : data_out = 24'b000000011011000001011011;
    16'b0000101001101011 : data_out = 24'b000000011011000011000111;
    16'b0000101001101100 : data_out = 24'b000000011011000100110011;
    16'b0000101001101101 : data_out = 24'b000000011011000110100000;
    16'b0000101001101110 : data_out = 24'b000000011011001000001100;
    16'b0000101001101111 : data_out = 24'b000000011011001001111001;
    16'b0000101001110000 : data_out = 24'b000000011011001011100101;
    16'b0000101001110001 : data_out = 24'b000000011011001101010010;
    16'b0000101001110010 : data_out = 24'b000000011011001110111111;
    16'b0000101001110011 : data_out = 24'b000000011011010000101100;
    16'b0000101001110100 : data_out = 24'b000000011011010010011001;
    16'b0000101001110101 : data_out = 24'b000000011011010100000110;
    16'b0000101001110110 : data_out = 24'b000000011011010101110100;
    16'b0000101001110111 : data_out = 24'b000000011011010111100001;
    16'b0000101001111000 : data_out = 24'b000000011011011001001111;
    16'b0000101001111001 : data_out = 24'b000000011011011010111100;
    16'b0000101001111010 : data_out = 24'b000000011011011100101010;
    16'b0000101001111011 : data_out = 24'b000000011011011110011000;
    16'b0000101001111100 : data_out = 24'b000000011011100000000110;
    16'b0000101001111101 : data_out = 24'b000000011011100001110100;
    16'b0000101001111110 : data_out = 24'b000000011011100011100010;
    16'b0000101001111111 : data_out = 24'b000000011011100101010000;
    16'b0000101010000000 : data_out = 24'b000000011011100110111111;
    16'b0000101010000001 : data_out = 24'b000000011011101000101101;
    16'b0000101010000010 : data_out = 24'b000000011011101010011100;
    16'b0000101010000011 : data_out = 24'b000000011011101100001010;
    16'b0000101010000100 : data_out = 24'b000000011011101101111001;
    16'b0000101010000101 : data_out = 24'b000000011011101111101000;
    16'b0000101010000110 : data_out = 24'b000000011011110001010111;
    16'b0000101010000111 : data_out = 24'b000000011011110011000110;
    16'b0000101010001000 : data_out = 24'b000000011011110100110110;
    16'b0000101010001001 : data_out = 24'b000000011011110110100101;
    16'b0000101010001010 : data_out = 24'b000000011011111000010100;
    16'b0000101010001011 : data_out = 24'b000000011011111010000100;
    16'b0000101010001100 : data_out = 24'b000000011011111011110100;
    16'b0000101010001101 : data_out = 24'b000000011011111101100011;
    16'b0000101010001110 : data_out = 24'b000000011011111111010011;
    16'b0000101010001111 : data_out = 24'b000000011100000001000011;
    16'b0000101010010000 : data_out = 24'b000000011100000010110011;
    16'b0000101010010001 : data_out = 24'b000000011100000100100100;
    16'b0000101010010010 : data_out = 24'b000000011100000110010100;
    16'b0000101010010011 : data_out = 24'b000000011100001000000100;
    16'b0000101010010100 : data_out = 24'b000000011100001001110101;
    16'b0000101010010101 : data_out = 24'b000000011100001011100110;
    16'b0000101010010110 : data_out = 24'b000000011100001101010110;
    16'b0000101010010111 : data_out = 24'b000000011100001111000111;
    16'b0000101010011000 : data_out = 24'b000000011100010000111000;
    16'b0000101010011001 : data_out = 24'b000000011100010010101001;
    16'b0000101010011010 : data_out = 24'b000000011100010100011011;
    16'b0000101010011011 : data_out = 24'b000000011100010110001100;
    16'b0000101010011100 : data_out = 24'b000000011100010111111101;
    16'b0000101010011101 : data_out = 24'b000000011100011001101111;
    16'b0000101010011110 : data_out = 24'b000000011100011011100001;
    16'b0000101010011111 : data_out = 24'b000000011100011101010010;
    16'b0000101010100000 : data_out = 24'b000000011100011111000100;
    16'b0000101010100001 : data_out = 24'b000000011100100000110110;
    16'b0000101010100010 : data_out = 24'b000000011100100010101000;
    16'b0000101010100011 : data_out = 24'b000000011100100100011011;
    16'b0000101010100100 : data_out = 24'b000000011100100110001101;
    16'b0000101010100101 : data_out = 24'b000000011100100111111111;
    16'b0000101010100110 : data_out = 24'b000000011100101001110010;
    16'b0000101010100111 : data_out = 24'b000000011100101011100101;
    16'b0000101010101000 : data_out = 24'b000000011100101101010111;
    16'b0000101010101001 : data_out = 24'b000000011100101111001010;
    16'b0000101010101010 : data_out = 24'b000000011100110000111101;
    16'b0000101010101011 : data_out = 24'b000000011100110010110000;
    16'b0000101010101100 : data_out = 24'b000000011100110100100100;
    16'b0000101010101101 : data_out = 24'b000000011100110110010111;
    16'b0000101010101110 : data_out = 24'b000000011100111000001010;
    16'b0000101010101111 : data_out = 24'b000000011100111001111110;
    16'b0000101010110000 : data_out = 24'b000000011100111011110010;
    16'b0000101010110001 : data_out = 24'b000000011100111101100110;
    16'b0000101010110010 : data_out = 24'b000000011100111111011001;
    16'b0000101010110011 : data_out = 24'b000000011101000001001101;
    16'b0000101010110100 : data_out = 24'b000000011101000011000010;
    16'b0000101010110101 : data_out = 24'b000000011101000100110110;
    16'b0000101010110110 : data_out = 24'b000000011101000110101010;
    16'b0000101010110111 : data_out = 24'b000000011101001000011111;
    16'b0000101010111000 : data_out = 24'b000000011101001010010011;
    16'b0000101010111001 : data_out = 24'b000000011101001100001000;
    16'b0000101010111010 : data_out = 24'b000000011101001101111101;
    16'b0000101010111011 : data_out = 24'b000000011101001111110010;
    16'b0000101010111100 : data_out = 24'b000000011101010001100111;
    16'b0000101010111101 : data_out = 24'b000000011101010011011100;
    16'b0000101010111110 : data_out = 24'b000000011101010101010001;
    16'b0000101010111111 : data_out = 24'b000000011101010111000111;
    16'b0000101011000000 : data_out = 24'b000000011101011000111100;
    16'b0000101011000001 : data_out = 24'b000000011101011010110010;
    16'b0000101011000010 : data_out = 24'b000000011101011100100111;
    16'b0000101011000011 : data_out = 24'b000000011101011110011101;
    16'b0000101011000100 : data_out = 24'b000000011101100000010011;
    16'b0000101011000101 : data_out = 24'b000000011101100010001001;
    16'b0000101011000110 : data_out = 24'b000000011101100011111111;
    16'b0000101011000111 : data_out = 24'b000000011101100101110110;
    16'b0000101011001000 : data_out = 24'b000000011101100111101100;
    16'b0000101011001001 : data_out = 24'b000000011101101001100011;
    16'b0000101011001010 : data_out = 24'b000000011101101011011001;
    16'b0000101011001011 : data_out = 24'b000000011101101101010000;
    16'b0000101011001100 : data_out = 24'b000000011101101111000111;
    16'b0000101011001101 : data_out = 24'b000000011101110000111110;
    16'b0000101011001110 : data_out = 24'b000000011101110010110101;
    16'b0000101011001111 : data_out = 24'b000000011101110100101100;
    16'b0000101011010000 : data_out = 24'b000000011101110110100100;
    16'b0000101011010001 : data_out = 24'b000000011101111000011011;
    16'b0000101011010010 : data_out = 24'b000000011101111010010011;
    16'b0000101011010011 : data_out = 24'b000000011101111100001011;
    16'b0000101011010100 : data_out = 24'b000000011101111110000010;
    16'b0000101011010101 : data_out = 24'b000000011101111111111010;
    16'b0000101011010110 : data_out = 24'b000000011110000001110010;
    16'b0000101011010111 : data_out = 24'b000000011110000011101011;
    16'b0000101011011000 : data_out = 24'b000000011110000101100011;
    16'b0000101011011001 : data_out = 24'b000000011110000111011011;
    16'b0000101011011010 : data_out = 24'b000000011110001001010100;
    16'b0000101011011011 : data_out = 24'b000000011110001011001100;
    16'b0000101011011100 : data_out = 24'b000000011110001101000101;
    16'b0000101011011101 : data_out = 24'b000000011110001110111110;
    16'b0000101011011110 : data_out = 24'b000000011110010000110111;
    16'b0000101011011111 : data_out = 24'b000000011110010010110000;
    16'b0000101011100000 : data_out = 24'b000000011110010100101001;
    16'b0000101011100001 : data_out = 24'b000000011110010110100011;
    16'b0000101011100010 : data_out = 24'b000000011110011000011100;
    16'b0000101011100011 : data_out = 24'b000000011110011010010110;
    16'b0000101011100100 : data_out = 24'b000000011110011100001111;
    16'b0000101011100101 : data_out = 24'b000000011110011110001001;
    16'b0000101011100110 : data_out = 24'b000000011110100000000011;
    16'b0000101011100111 : data_out = 24'b000000011110100001111101;
    16'b0000101011101000 : data_out = 24'b000000011110100011110111;
    16'b0000101011101001 : data_out = 24'b000000011110100101110010;
    16'b0000101011101010 : data_out = 24'b000000011110100111101100;
    16'b0000101011101011 : data_out = 24'b000000011110101001100111;
    16'b0000101011101100 : data_out = 24'b000000011110101011100001;
    16'b0000101011101101 : data_out = 24'b000000011110101101011100;
    16'b0000101011101110 : data_out = 24'b000000011110101111010111;
    16'b0000101011101111 : data_out = 24'b000000011110110001010010;
    16'b0000101011110000 : data_out = 24'b000000011110110011001101;
    16'b0000101011110001 : data_out = 24'b000000011110110101001001;
    16'b0000101011110010 : data_out = 24'b000000011110110111000100;
    16'b0000101011110011 : data_out = 24'b000000011110111000111111;
    16'b0000101011110100 : data_out = 24'b000000011110111010111011;
    16'b0000101011110101 : data_out = 24'b000000011110111100110111;
    16'b0000101011110110 : data_out = 24'b000000011110111110110011;
    16'b0000101011110111 : data_out = 24'b000000011111000000101111;
    16'b0000101011111000 : data_out = 24'b000000011111000010101011;
    16'b0000101011111001 : data_out = 24'b000000011111000100100111;
    16'b0000101011111010 : data_out = 24'b000000011111000110100011;
    16'b0000101011111011 : data_out = 24'b000000011111001000100000;
    16'b0000101011111100 : data_out = 24'b000000011111001010011100;
    16'b0000101011111101 : data_out = 24'b000000011111001100011001;
    16'b0000101011111110 : data_out = 24'b000000011111001110010110;
    16'b0000101011111111 : data_out = 24'b000000011111010000010011;
    16'b0000101100000000 : data_out = 24'b000000011111010010010000;
    16'b0000101100000001 : data_out = 24'b000000011111010100001101;
    16'b0000101100000010 : data_out = 24'b000000011111010110001010;
    16'b0000101100000011 : data_out = 24'b000000011111011000001000;
    16'b0000101100000100 : data_out = 24'b000000011111011010000101;
    16'b0000101100000101 : data_out = 24'b000000011111011100000011;
    16'b0000101100000110 : data_out = 24'b000000011111011110000001;
    16'b0000101100000111 : data_out = 24'b000000011111011111111111;
    16'b0000101100001000 : data_out = 24'b000000011111100001111101;
    16'b0000101100001001 : data_out = 24'b000000011111100011111011;
    16'b0000101100001010 : data_out = 24'b000000011111100101111001;
    16'b0000101100001011 : data_out = 24'b000000011111100111111000;
    16'b0000101100001100 : data_out = 24'b000000011111101001110110;
    16'b0000101100001101 : data_out = 24'b000000011111101011110101;
    16'b0000101100001110 : data_out = 24'b000000011111101101110100;
    16'b0000101100001111 : data_out = 24'b000000011111101111110011;
    16'b0000101100010000 : data_out = 24'b000000011111110001110010;
    16'b0000101100010001 : data_out = 24'b000000011111110011110001;
    16'b0000101100010010 : data_out = 24'b000000011111110101110000;
    16'b0000101100010011 : data_out = 24'b000000011111110111110000;
    16'b0000101100010100 : data_out = 24'b000000011111111001101111;
    16'b0000101100010101 : data_out = 24'b000000011111111011101111;
    16'b0000101100010110 : data_out = 24'b000000011111111101101111;
    16'b0000101100010111 : data_out = 24'b000000011111111111101111;
    16'b0000101100011000 : data_out = 24'b000000100000000001101111;
    16'b0000101100011001 : data_out = 24'b000000100000000011101111;
    16'b0000101100011010 : data_out = 24'b000000100000000101101111;
    16'b0000101100011011 : data_out = 24'b000000100000000111110000;
    16'b0000101100011100 : data_out = 24'b000000100000001001110000;
    16'b0000101100011101 : data_out = 24'b000000100000001011110001;
    16'b0000101100011110 : data_out = 24'b000000100000001101110010;
    16'b0000101100011111 : data_out = 24'b000000100000001111110011;
    16'b0000101100100000 : data_out = 24'b000000100000010001110100;
    16'b0000101100100001 : data_out = 24'b000000100000010011110101;
    16'b0000101100100010 : data_out = 24'b000000100000010101110110;
    16'b0000101100100011 : data_out = 24'b000000100000010111111000;
    16'b0000101100100100 : data_out = 24'b000000100000011001111001;
    16'b0000101100100101 : data_out = 24'b000000100000011011111011;
    16'b0000101100100110 : data_out = 24'b000000100000011101111101;
    16'b0000101100100111 : data_out = 24'b000000100000011111111111;
    16'b0000101100101000 : data_out = 24'b000000100000100010000001;
    16'b0000101100101001 : data_out = 24'b000000100000100100000011;
    16'b0000101100101010 : data_out = 24'b000000100000100110000101;
    16'b0000101100101011 : data_out = 24'b000000100000101000001000;
    16'b0000101100101100 : data_out = 24'b000000100000101010001010;
    16'b0000101100101101 : data_out = 24'b000000100000101100001101;
    16'b0000101100101110 : data_out = 24'b000000100000101110010000;
    16'b0000101100101111 : data_out = 24'b000000100000110000010011;
    16'b0000101100110000 : data_out = 24'b000000100000110010010110;
    16'b0000101100110001 : data_out = 24'b000000100000110100011001;
    16'b0000101100110010 : data_out = 24'b000000100000110110011100;
    16'b0000101100110011 : data_out = 24'b000000100000111000100000;
    16'b0000101100110100 : data_out = 24'b000000100000111010100011;
    16'b0000101100110101 : data_out = 24'b000000100000111100100111;
    16'b0000101100110110 : data_out = 24'b000000100000111110101011;
    16'b0000101100110111 : data_out = 24'b000000100001000000101111;
    16'b0000101100111000 : data_out = 24'b000000100001000010110011;
    16'b0000101100111001 : data_out = 24'b000000100001000100110111;
    16'b0000101100111010 : data_out = 24'b000000100001000110111100;
    16'b0000101100111011 : data_out = 24'b000000100001001001000000;
    16'b0000101100111100 : data_out = 24'b000000100001001011000101;
    16'b0000101100111101 : data_out = 24'b000000100001001101001001;
    16'b0000101100111110 : data_out = 24'b000000100001001111001110;
    16'b0000101100111111 : data_out = 24'b000000100001010001010011;
    16'b0000101101000000 : data_out = 24'b000000100001010011011001;
    16'b0000101101000001 : data_out = 24'b000000100001010101011110;
    16'b0000101101000010 : data_out = 24'b000000100001010111100011;
    16'b0000101101000011 : data_out = 24'b000000100001011001101001;
    16'b0000101101000100 : data_out = 24'b000000100001011011101110;
    16'b0000101101000101 : data_out = 24'b000000100001011101110100;
    16'b0000101101000110 : data_out = 24'b000000100001011111111010;
    16'b0000101101000111 : data_out = 24'b000000100001100010000000;
    16'b0000101101001000 : data_out = 24'b000000100001100100000110;
    16'b0000101101001001 : data_out = 24'b000000100001100110001101;
    16'b0000101101001010 : data_out = 24'b000000100001101000010011;
    16'b0000101101001011 : data_out = 24'b000000100001101010011010;
    16'b0000101101001100 : data_out = 24'b000000100001101100100000;
    16'b0000101101001101 : data_out = 24'b000000100001101110100111;
    16'b0000101101001110 : data_out = 24'b000000100001110000101110;
    16'b0000101101001111 : data_out = 24'b000000100001110010110101;
    16'b0000101101010000 : data_out = 24'b000000100001110100111101;
    16'b0000101101010001 : data_out = 24'b000000100001110111000100;
    16'b0000101101010010 : data_out = 24'b000000100001111001001100;
    16'b0000101101010011 : data_out = 24'b000000100001111011010011;
    16'b0000101101010100 : data_out = 24'b000000100001111101011011;
    16'b0000101101010101 : data_out = 24'b000000100001111111100011;
    16'b0000101101010110 : data_out = 24'b000000100010000001101011;
    16'b0000101101010111 : data_out = 24'b000000100010000011110011;
    16'b0000101101011000 : data_out = 24'b000000100010000101111011;
    16'b0000101101011001 : data_out = 24'b000000100010001000000100;
    16'b0000101101011010 : data_out = 24'b000000100010001010001100;
    16'b0000101101011011 : data_out = 24'b000000100010001100010101;
    16'b0000101101011100 : data_out = 24'b000000100010001110011110;
    16'b0000101101011101 : data_out = 24'b000000100010010000100111;
    16'b0000101101011110 : data_out = 24'b000000100010010010110000;
    16'b0000101101011111 : data_out = 24'b000000100010010100111001;
    16'b0000101101100000 : data_out = 24'b000000100010010111000011;
    16'b0000101101100001 : data_out = 24'b000000100010011001001100;
    16'b0000101101100010 : data_out = 24'b000000100010011011010110;
    16'b0000101101100011 : data_out = 24'b000000100010011101100000;
    16'b0000101101100100 : data_out = 24'b000000100010011111101001;
    16'b0000101101100101 : data_out = 24'b000000100010100001110100;
    16'b0000101101100110 : data_out = 24'b000000100010100011111110;
    16'b0000101101100111 : data_out = 24'b000000100010100110001000;
    16'b0000101101101000 : data_out = 24'b000000100010101000010010;
    16'b0000101101101001 : data_out = 24'b000000100010101010011101;
    16'b0000101101101010 : data_out = 24'b000000100010101100101000;
    16'b0000101101101011 : data_out = 24'b000000100010101110110011;
    16'b0000101101101100 : data_out = 24'b000000100010110000111110;
    16'b0000101101101101 : data_out = 24'b000000100010110011001001;
    16'b0000101101101110 : data_out = 24'b000000100010110101010100;
    16'b0000101101101111 : data_out = 24'b000000100010110111011111;
    16'b0000101101110000 : data_out = 24'b000000100010111001101011;
    16'b0000101101110001 : data_out = 24'b000000100010111011110111;
    16'b0000101101110010 : data_out = 24'b000000100010111110000010;
    16'b0000101101110011 : data_out = 24'b000000100011000000001110;
    16'b0000101101110100 : data_out = 24'b000000100011000010011010;
    16'b0000101101110101 : data_out = 24'b000000100011000100100111;
    16'b0000101101110110 : data_out = 24'b000000100011000110110011;
    16'b0000101101110111 : data_out = 24'b000000100011001001000000;
    16'b0000101101111000 : data_out = 24'b000000100011001011001100;
    16'b0000101101111001 : data_out = 24'b000000100011001101011001;
    16'b0000101101111010 : data_out = 24'b000000100011001111100110;
    16'b0000101101111011 : data_out = 24'b000000100011010001110011;
    16'b0000101101111100 : data_out = 24'b000000100011010100000000;
    16'b0000101101111101 : data_out = 24'b000000100011010110001101;
    16'b0000101101111110 : data_out = 24'b000000100011011000011011;
    16'b0000101101111111 : data_out = 24'b000000100011011010101000;
    16'b0000101110000000 : data_out = 24'b000000100011011100110110;
    16'b0000101110000001 : data_out = 24'b000000100011011111000100;
    16'b0000101110000010 : data_out = 24'b000000100011100001010010;
    16'b0000101110000011 : data_out = 24'b000000100011100011100000;
    16'b0000101110000100 : data_out = 24'b000000100011100101101110;
    16'b0000101110000101 : data_out = 24'b000000100011100111111101;
    16'b0000101110000110 : data_out = 24'b000000100011101010001011;
    16'b0000101110000111 : data_out = 24'b000000100011101100011010;
    16'b0000101110001000 : data_out = 24'b000000100011101110101001;
    16'b0000101110001001 : data_out = 24'b000000100011110000111000;
    16'b0000101110001010 : data_out = 24'b000000100011110011000111;
    16'b0000101110001011 : data_out = 24'b000000100011110101010110;
    16'b0000101110001100 : data_out = 24'b000000100011110111100110;
    16'b0000101110001101 : data_out = 24'b000000100011111001110101;
    16'b0000101110001110 : data_out = 24'b000000100011111100000101;
    16'b0000101110001111 : data_out = 24'b000000100011111110010101;
    16'b0000101110010000 : data_out = 24'b000000100100000000100101;
    16'b0000101110010001 : data_out = 24'b000000100100000010110101;
    16'b0000101110010010 : data_out = 24'b000000100100000101000101;
    16'b0000101110010011 : data_out = 24'b000000100100000111010110;
    16'b0000101110010100 : data_out = 24'b000000100100001001100110;
    16'b0000101110010101 : data_out = 24'b000000100100001011110111;
    16'b0000101110010110 : data_out = 24'b000000100100001110001000;
    16'b0000101110010111 : data_out = 24'b000000100100010000011001;
    16'b0000101110011000 : data_out = 24'b000000100100010010101010;
    16'b0000101110011001 : data_out = 24'b000000100100010100111011;
    16'b0000101110011010 : data_out = 24'b000000100100010111001100;
    16'b0000101110011011 : data_out = 24'b000000100100011001011110;
    16'b0000101110011100 : data_out = 24'b000000100100011011101111;
    16'b0000101110011101 : data_out = 24'b000000100100011110000001;
    16'b0000101110011110 : data_out = 24'b000000100100100000010011;
    16'b0000101110011111 : data_out = 24'b000000100100100010100101;
    16'b0000101110100000 : data_out = 24'b000000100100100100111000;
    16'b0000101110100001 : data_out = 24'b000000100100100111001010;
    16'b0000101110100010 : data_out = 24'b000000100100101001011100;
    16'b0000101110100011 : data_out = 24'b000000100100101011101111;
    16'b0000101110100100 : data_out = 24'b000000100100101110000010;
    16'b0000101110100101 : data_out = 24'b000000100100110000010101;
    16'b0000101110100110 : data_out = 24'b000000100100110010101000;
    16'b0000101110100111 : data_out = 24'b000000100100110100111011;
    16'b0000101110101000 : data_out = 24'b000000100100110111001111;
    16'b0000101110101001 : data_out = 24'b000000100100111001100010;
    16'b0000101110101010 : data_out = 24'b000000100100111011110110;
    16'b0000101110101011 : data_out = 24'b000000100100111110001010;
    16'b0000101110101100 : data_out = 24'b000000100101000000011110;
    16'b0000101110101101 : data_out = 24'b000000100101000010110010;
    16'b0000101110101110 : data_out = 24'b000000100101000101000110;
    16'b0000101110101111 : data_out = 24'b000000100101000111011010;
    16'b0000101110110000 : data_out = 24'b000000100101001001101111;
    16'b0000101110110001 : data_out = 24'b000000100101001100000011;
    16'b0000101110110010 : data_out = 24'b000000100101001110011000;
    16'b0000101110110011 : data_out = 24'b000000100101010000101101;
    16'b0000101110110100 : data_out = 24'b000000100101010011000010;
    16'b0000101110110101 : data_out = 24'b000000100101010101011000;
    16'b0000101110110110 : data_out = 24'b000000100101010111101101;
    16'b0000101110110111 : data_out = 24'b000000100101011010000011;
    16'b0000101110111000 : data_out = 24'b000000100101011100011000;
    16'b0000101110111001 : data_out = 24'b000000100101011110101110;
    16'b0000101110111010 : data_out = 24'b000000100101100001000100;
    16'b0000101110111011 : data_out = 24'b000000100101100011011010;
    16'b0000101110111100 : data_out = 24'b000000100101100101110001;
    16'b0000101110111101 : data_out = 24'b000000100101101000000111;
    16'b0000101110111110 : data_out = 24'b000000100101101010011110;
    16'b0000101110111111 : data_out = 24'b000000100101101100110100;
    16'b0000101111000000 : data_out = 24'b000000100101101111001011;
    16'b0000101111000001 : data_out = 24'b000000100101110001100010;
    16'b0000101111000010 : data_out = 24'b000000100101110011111001;
    16'b0000101111000011 : data_out = 24'b000000100101110110010001;
    16'b0000101111000100 : data_out = 24'b000000100101111000101000;
    16'b0000101111000101 : data_out = 24'b000000100101111011000000;
    16'b0000101111000110 : data_out = 24'b000000100101111101011000;
    16'b0000101111000111 : data_out = 24'b000000100101111111101111;
    16'b0000101111001000 : data_out = 24'b000000100110000010001000;
    16'b0000101111001001 : data_out = 24'b000000100110000100100000;
    16'b0000101111001010 : data_out = 24'b000000100110000110111000;
    16'b0000101111001011 : data_out = 24'b000000100110001001010001;
    16'b0000101111001100 : data_out = 24'b000000100110001011101001;
    16'b0000101111001101 : data_out = 24'b000000100110001110000010;
    16'b0000101111001110 : data_out = 24'b000000100110010000011011;
    16'b0000101111001111 : data_out = 24'b000000100110010010110100;
    16'b0000101111010000 : data_out = 24'b000000100110010101001101;
    16'b0000101111010001 : data_out = 24'b000000100110010111100111;
    16'b0000101111010010 : data_out = 24'b000000100110011010000000;
    16'b0000101111010011 : data_out = 24'b000000100110011100011010;
    16'b0000101111010100 : data_out = 24'b000000100110011110110100;
    16'b0000101111010101 : data_out = 24'b000000100110100001001110;
    16'b0000101111010110 : data_out = 24'b000000100110100011101000;
    16'b0000101111010111 : data_out = 24'b000000100110100110000010;
    16'b0000101111011000 : data_out = 24'b000000100110101000011101;
    16'b0000101111011001 : data_out = 24'b000000100110101010110111;
    16'b0000101111011010 : data_out = 24'b000000100110101101010010;
    16'b0000101111011011 : data_out = 24'b000000100110101111101101;
    16'b0000101111011100 : data_out = 24'b000000100110110010001000;
    16'b0000101111011101 : data_out = 24'b000000100110110100100011;
    16'b0000101111011110 : data_out = 24'b000000100110110110111111;
    16'b0000101111011111 : data_out = 24'b000000100110111001011010;
    16'b0000101111100000 : data_out = 24'b000000100110111011110110;
    16'b0000101111100001 : data_out = 24'b000000100110111110010010;
    16'b0000101111100010 : data_out = 24'b000000100111000000101110;
    16'b0000101111100011 : data_out = 24'b000000100111000011001010;
    16'b0000101111100100 : data_out = 24'b000000100111000101100110;
    16'b0000101111100101 : data_out = 24'b000000100111001000000010;
    16'b0000101111100110 : data_out = 24'b000000100111001010011111;
    16'b0000101111100111 : data_out = 24'b000000100111001100111100;
    16'b0000101111101000 : data_out = 24'b000000100111001111011001;
    16'b0000101111101001 : data_out = 24'b000000100111010001110110;
    16'b0000101111101010 : data_out = 24'b000000100111010100010011;
    16'b0000101111101011 : data_out = 24'b000000100111010110110000;
    16'b0000101111101100 : data_out = 24'b000000100111011001001110;
    16'b0000101111101101 : data_out = 24'b000000100111011011101011;
    16'b0000101111101110 : data_out = 24'b000000100111011110001001;
    16'b0000101111101111 : data_out = 24'b000000100111100000100111;
    16'b0000101111110000 : data_out = 24'b000000100111100011000101;
    16'b0000101111110001 : data_out = 24'b000000100111100101100100;
    16'b0000101111110010 : data_out = 24'b000000100111101000000010;
    16'b0000101111110011 : data_out = 24'b000000100111101010100001;
    16'b0000101111110100 : data_out = 24'b000000100111101100111111;
    16'b0000101111110101 : data_out = 24'b000000100111101111011110;
    16'b0000101111110110 : data_out = 24'b000000100111110001111101;
    16'b0000101111110111 : data_out = 24'b000000100111110100011100;
    16'b0000101111111000 : data_out = 24'b000000100111110110111100;
    16'b0000101111111001 : data_out = 24'b000000100111111001011011;
    16'b0000101111111010 : data_out = 24'b000000100111111011111011;
    16'b0000101111111011 : data_out = 24'b000000100111111110011011;
    16'b0000101111111100 : data_out = 24'b000000101000000000111011;
    16'b0000101111111101 : data_out = 24'b000000101000000011011011;
    16'b0000101111111110 : data_out = 24'b000000101000000101111011;
    16'b0000101111111111 : data_out = 24'b000000101000001000011100;
    16'b0000110000000000 : data_out = 24'b000000101000001010111100;
    16'b0000110000000001 : data_out = 24'b000000101000001101011101;
    16'b0000110000000010 : data_out = 24'b000000101000001111111110;
    16'b0000110000000011 : data_out = 24'b000000101000010010011111;
    16'b0000110000000100 : data_out = 24'b000000101000010101000000;
    16'b0000110000000101 : data_out = 24'b000000101000010111100010;
    16'b0000110000000110 : data_out = 24'b000000101000011010000011;
    16'b0000110000000111 : data_out = 24'b000000101000011100100101;
    16'b0000110000001000 : data_out = 24'b000000101000011111000111;
    16'b0000110000001001 : data_out = 24'b000000101000100001101001;
    16'b0000110000001010 : data_out = 24'b000000101000100100001011;
    16'b0000110000001011 : data_out = 24'b000000101000100110101101;
    16'b0000110000001100 : data_out = 24'b000000101000101001010000;
    16'b0000110000001101 : data_out = 24'b000000101000101011110010;
    16'b0000110000001110 : data_out = 24'b000000101000101110010101;
    16'b0000110000001111 : data_out = 24'b000000101000110000111000;
    16'b0000110000010000 : data_out = 24'b000000101000110011011011;
    16'b0000110000010001 : data_out = 24'b000000101000110101111111;
    16'b0000110000010010 : data_out = 24'b000000101000111000100010;
    16'b0000110000010011 : data_out = 24'b000000101000111011000110;
    16'b0000110000010100 : data_out = 24'b000000101000111101101001;
    16'b0000110000010101 : data_out = 24'b000000101001000000001101;
    16'b0000110000010110 : data_out = 24'b000000101001000010110010;
    16'b0000110000010111 : data_out = 24'b000000101001000101010110;
    16'b0000110000011000 : data_out = 24'b000000101001000111111010;
    16'b0000110000011001 : data_out = 24'b000000101001001010011111;
    16'b0000110000011010 : data_out = 24'b000000101001001101000100;
    16'b0000110000011011 : data_out = 24'b000000101001001111101000;
    16'b0000110000011100 : data_out = 24'b000000101001010010001101;
    16'b0000110000011101 : data_out = 24'b000000101001010100110011;
    16'b0000110000011110 : data_out = 24'b000000101001010111011000;
    16'b0000110000011111 : data_out = 24'b000000101001011001111110;
    16'b0000110000100000 : data_out = 24'b000000101001011100100011;
    16'b0000110000100001 : data_out = 24'b000000101001011111001001;
    16'b0000110000100010 : data_out = 24'b000000101001100001101111;
    16'b0000110000100011 : data_out = 24'b000000101001100100010101;
    16'b0000110000100100 : data_out = 24'b000000101001100110111100;
    16'b0000110000100101 : data_out = 24'b000000101001101001100010;
    16'b0000110000100110 : data_out = 24'b000000101001101100001001;
    16'b0000110000100111 : data_out = 24'b000000101001101110110000;
    16'b0000110000101000 : data_out = 24'b000000101001110001010111;
    16'b0000110000101001 : data_out = 24'b000000101001110011111110;
    16'b0000110000101010 : data_out = 24'b000000101001110110100101;
    16'b0000110000101011 : data_out = 24'b000000101001111001001101;
    16'b0000110000101100 : data_out = 24'b000000101001111011110100;
    16'b0000110000101101 : data_out = 24'b000000101001111110011100;
    16'b0000110000101110 : data_out = 24'b000000101010000001000100;
    16'b0000110000101111 : data_out = 24'b000000101010000011101100;
    16'b0000110000110000 : data_out = 24'b000000101010000110010101;
    16'b0000110000110001 : data_out = 24'b000000101010001000111101;
    16'b0000110000110010 : data_out = 24'b000000101010001011100110;
    16'b0000110000110011 : data_out = 24'b000000101010001110001111;
    16'b0000110000110100 : data_out = 24'b000000101010010000111000;
    16'b0000110000110101 : data_out = 24'b000000101010010011100001;
    16'b0000110000110110 : data_out = 24'b000000101010010110001010;
    16'b0000110000110111 : data_out = 24'b000000101010011000110100;
    16'b0000110000111000 : data_out = 24'b000000101010011011011101;
    16'b0000110000111001 : data_out = 24'b000000101010011110000111;
    16'b0000110000111010 : data_out = 24'b000000101010100000110001;
    16'b0000110000111011 : data_out = 24'b000000101010100011011011;
    16'b0000110000111100 : data_out = 24'b000000101010100110000101;
    16'b0000110000111101 : data_out = 24'b000000101010101000110000;
    16'b0000110000111110 : data_out = 24'b000000101010101011011010;
    16'b0000110000111111 : data_out = 24'b000000101010101110000101;
    16'b0000110001000000 : data_out = 24'b000000101010110000110000;
    16'b0000110001000001 : data_out = 24'b000000101010110011011011;
    16'b0000110001000010 : data_out = 24'b000000101010110110000111;
    16'b0000110001000011 : data_out = 24'b000000101010111000110010;
    16'b0000110001000100 : data_out = 24'b000000101010111011011110;
    16'b0000110001000101 : data_out = 24'b000000101010111110001010;
    16'b0000110001000110 : data_out = 24'b000000101011000000110101;
    16'b0000110001000111 : data_out = 24'b000000101011000011100010;
    16'b0000110001001000 : data_out = 24'b000000101011000110001110;
    16'b0000110001001001 : data_out = 24'b000000101011001000111010;
    16'b0000110001001010 : data_out = 24'b000000101011001011100111;
    16'b0000110001001011 : data_out = 24'b000000101011001110010100;
    16'b0000110001001100 : data_out = 24'b000000101011010001000001;
    16'b0000110001001101 : data_out = 24'b000000101011010011101110;
    16'b0000110001001110 : data_out = 24'b000000101011010110011011;
    16'b0000110001001111 : data_out = 24'b000000101011011001001001;
    16'b0000110001010000 : data_out = 24'b000000101011011011110110;
    16'b0000110001010001 : data_out = 24'b000000101011011110100100;
    16'b0000110001010010 : data_out = 24'b000000101011100001010010;
    16'b0000110001010011 : data_out = 24'b000000101011100100000000;
    16'b0000110001010100 : data_out = 24'b000000101011100110101111;
    16'b0000110001010101 : data_out = 24'b000000101011101001011101;
    16'b0000110001010110 : data_out = 24'b000000101011101100001100;
    16'b0000110001010111 : data_out = 24'b000000101011101110111011;
    16'b0000110001011000 : data_out = 24'b000000101011110001101010;
    16'b0000110001011001 : data_out = 24'b000000101011110100011001;
    16'b0000110001011010 : data_out = 24'b000000101011110111001000;
    16'b0000110001011011 : data_out = 24'b000000101011111001111000;
    16'b0000110001011100 : data_out = 24'b000000101011111100101000;
    16'b0000110001011101 : data_out = 24'b000000101011111111010111;
    16'b0000110001011110 : data_out = 24'b000000101100000010001000;
    16'b0000110001011111 : data_out = 24'b000000101100000100111000;
    16'b0000110001100000 : data_out = 24'b000000101100000111101000;
    16'b0000110001100001 : data_out = 24'b000000101100001010011001;
    16'b0000110001100010 : data_out = 24'b000000101100001101001001;
    16'b0000110001100011 : data_out = 24'b000000101100001111111010;
    16'b0000110001100100 : data_out = 24'b000000101100010010101011;
    16'b0000110001100101 : data_out = 24'b000000101100010101011101;
    16'b0000110001100110 : data_out = 24'b000000101100011000001110;
    16'b0000110001100111 : data_out = 24'b000000101100011011000000;
    16'b0000110001101000 : data_out = 24'b000000101100011101110001;
    16'b0000110001101001 : data_out = 24'b000000101100100000100011;
    16'b0000110001101010 : data_out = 24'b000000101100100011010110;
    16'b0000110001101011 : data_out = 24'b000000101100100110001000;
    16'b0000110001101100 : data_out = 24'b000000101100101000111010;
    16'b0000110001101101 : data_out = 24'b000000101100101011101101;
    16'b0000110001101110 : data_out = 24'b000000101100101110100000;
    16'b0000110001101111 : data_out = 24'b000000101100110001010011;
    16'b0000110001110000 : data_out = 24'b000000101100110100000110;
    16'b0000110001110001 : data_out = 24'b000000101100110110111001;
    16'b0000110001110010 : data_out = 24'b000000101100111001101101;
    16'b0000110001110011 : data_out = 24'b000000101100111100100000;
    16'b0000110001110100 : data_out = 24'b000000101100111111010100;
    16'b0000110001110101 : data_out = 24'b000000101101000010001000;
    16'b0000110001110110 : data_out = 24'b000000101101000100111101;
    16'b0000110001110111 : data_out = 24'b000000101101000111110001;
    16'b0000110001111000 : data_out = 24'b000000101101001010100110;
    16'b0000110001111001 : data_out = 24'b000000101101001101011010;
    16'b0000110001111010 : data_out = 24'b000000101101010000001111;
    16'b0000110001111011 : data_out = 24'b000000101101010011000100;
    16'b0000110001111100 : data_out = 24'b000000101101010101111010;
    16'b0000110001111101 : data_out = 24'b000000101101011000101111;
    16'b0000110001111110 : data_out = 24'b000000101101011011100101;
    16'b0000110001111111 : data_out = 24'b000000101101011110011011;
    16'b0000110010000000 : data_out = 24'b000000101101100001010001;
    16'b0000110010000001 : data_out = 24'b000000101101100100000111;
    16'b0000110010000010 : data_out = 24'b000000101101100110111101;
    16'b0000110010000011 : data_out = 24'b000000101101101001110100;
    16'b0000110010000100 : data_out = 24'b000000101101101100101010;
    16'b0000110010000101 : data_out = 24'b000000101101101111100001;
    16'b0000110010000110 : data_out = 24'b000000101101110010011000;
    16'b0000110010000111 : data_out = 24'b000000101101110101001111;
    16'b0000110010001000 : data_out = 24'b000000101101111000000111;
    16'b0000110010001001 : data_out = 24'b000000101101111010111110;
    16'b0000110010001010 : data_out = 24'b000000101101111101110110;
    16'b0000110010001011 : data_out = 24'b000000101110000000101110;
    16'b0000110010001100 : data_out = 24'b000000101110000011100110;
    16'b0000110010001101 : data_out = 24'b000000101110000110011111;
    16'b0000110010001110 : data_out = 24'b000000101110001001010111;
    16'b0000110010001111 : data_out = 24'b000000101110001100010000;
    16'b0000110010010000 : data_out = 24'b000000101110001111001001;
    16'b0000110010010001 : data_out = 24'b000000101110010010000010;
    16'b0000110010010010 : data_out = 24'b000000101110010100111011;
    16'b0000110010010011 : data_out = 24'b000000101110010111110100;
    16'b0000110010010100 : data_out = 24'b000000101110011010101110;
    16'b0000110010010101 : data_out = 24'b000000101110011101101000;
    16'b0000110010010110 : data_out = 24'b000000101110100000100010;
    16'b0000110010010111 : data_out = 24'b000000101110100011011100;
    16'b0000110010011000 : data_out = 24'b000000101110100110010110;
    16'b0000110010011001 : data_out = 24'b000000101110101001010001;
    16'b0000110010011010 : data_out = 24'b000000101110101100001011;
    16'b0000110010011011 : data_out = 24'b000000101110101111000110;
    16'b0000110010011100 : data_out = 24'b000000101110110010000001;
    16'b0000110010011101 : data_out = 24'b000000101110110100111100;
    16'b0000110010011110 : data_out = 24'b000000101110110111111000;
    16'b0000110010011111 : data_out = 24'b000000101110111010110011;
    16'b0000110010100000 : data_out = 24'b000000101110111101101111;
    16'b0000110010100001 : data_out = 24'b000000101111000000101011;
    16'b0000110010100010 : data_out = 24'b000000101111000011100111;
    16'b0000110010100011 : data_out = 24'b000000101111000110100011;
    16'b0000110010100100 : data_out = 24'b000000101111001001100000;
    16'b0000110010100101 : data_out = 24'b000000101111001100011101;
    16'b0000110010100110 : data_out = 24'b000000101111001111011010;
    16'b0000110010100111 : data_out = 24'b000000101111010010010111;
    16'b0000110010101000 : data_out = 24'b000000101111010101010100;
    16'b0000110010101001 : data_out = 24'b000000101111011000010001;
    16'b0000110010101010 : data_out = 24'b000000101111011011001111;
    16'b0000110010101011 : data_out = 24'b000000101111011110001101;
    16'b0000110010101100 : data_out = 24'b000000101111100001001011;
    16'b0000110010101101 : data_out = 24'b000000101111100100001001;
    16'b0000110010101110 : data_out = 24'b000000101111100111000111;
    16'b0000110010101111 : data_out = 24'b000000101111101010000110;
    16'b0000110010110000 : data_out = 24'b000000101111101101000100;
    16'b0000110010110001 : data_out = 24'b000000101111110000000011;
    16'b0000110010110010 : data_out = 24'b000000101111110011000010;
    16'b0000110010110011 : data_out = 24'b000000101111110110000010;
    16'b0000110010110100 : data_out = 24'b000000101111111001000001;
    16'b0000110010110101 : data_out = 24'b000000101111111100000001;
    16'b0000110010110110 : data_out = 24'b000000101111111111000001;
    16'b0000110010110111 : data_out = 24'b000000110000000010000001;
    16'b0000110010111000 : data_out = 24'b000000110000000101000001;
    16'b0000110010111001 : data_out = 24'b000000110000001000000001;
    16'b0000110010111010 : data_out = 24'b000000110000001011000010;
    16'b0000110010111011 : data_out = 24'b000000110000001110000011;
    16'b0000110010111100 : data_out = 24'b000000110000010001000100;
    16'b0000110010111101 : data_out = 24'b000000110000010100000101;
    16'b0000110010111110 : data_out = 24'b000000110000010111000110;
    16'b0000110010111111 : data_out = 24'b000000110000011010001000;
    16'b0000110011000000 : data_out = 24'b000000110000011101001001;
    16'b0000110011000001 : data_out = 24'b000000110000100000001011;
    16'b0000110011000010 : data_out = 24'b000000110000100011001110;
    16'b0000110011000011 : data_out = 24'b000000110000100110010000;
    16'b0000110011000100 : data_out = 24'b000000110000101001010010;
    16'b0000110011000101 : data_out = 24'b000000110000101100010101;
    16'b0000110011000110 : data_out = 24'b000000110000101111011000;
    16'b0000110011000111 : data_out = 24'b000000110000110010011011;
    16'b0000110011001000 : data_out = 24'b000000110000110101011110;
    16'b0000110011001001 : data_out = 24'b000000110000111000100010;
    16'b0000110011001010 : data_out = 24'b000000110000111011100101;
    16'b0000110011001011 : data_out = 24'b000000110000111110101001;
    16'b0000110011001100 : data_out = 24'b000000110001000001101101;
    16'b0000110011001101 : data_out = 24'b000000110001000100110001;
    16'b0000110011001110 : data_out = 24'b000000110001000111110110;
    16'b0000110011001111 : data_out = 24'b000000110001001010111010;
    16'b0000110011010000 : data_out = 24'b000000110001001101111111;
    16'b0000110011010001 : data_out = 24'b000000110001010001000100;
    16'b0000110011010010 : data_out = 24'b000000110001010100001001;
    16'b0000110011010011 : data_out = 24'b000000110001010111001110;
    16'b0000110011010100 : data_out = 24'b000000110001011010010100;
    16'b0000110011010101 : data_out = 24'b000000110001011101011010;
    16'b0000110011010110 : data_out = 24'b000000110001100000100000;
    16'b0000110011010111 : data_out = 24'b000000110001100011100110;
    16'b0000110011011000 : data_out = 24'b000000110001100110101100;
    16'b0000110011011001 : data_out = 24'b000000110001101001110011;
    16'b0000110011011010 : data_out = 24'b000000110001101100111001;
    16'b0000110011011011 : data_out = 24'b000000110001110000000000;
    16'b0000110011011100 : data_out = 24'b000000110001110011000111;
    16'b0000110011011101 : data_out = 24'b000000110001110110001111;
    16'b0000110011011110 : data_out = 24'b000000110001111001010110;
    16'b0000110011011111 : data_out = 24'b000000110001111100011110;
    16'b0000110011100000 : data_out = 24'b000000110001111111100110;
    16'b0000110011100001 : data_out = 24'b000000110010000010101110;
    16'b0000110011100010 : data_out = 24'b000000110010000101110110;
    16'b0000110011100011 : data_out = 24'b000000110010001000111111;
    16'b0000110011100100 : data_out = 24'b000000110010001100000111;
    16'b0000110011100101 : data_out = 24'b000000110010001111010000;
    16'b0000110011100110 : data_out = 24'b000000110010010010011001;
    16'b0000110011100111 : data_out = 24'b000000110010010101100010;
    16'b0000110011101000 : data_out = 24'b000000110010011000101100;
    16'b0000110011101001 : data_out = 24'b000000110010011011110101;
    16'b0000110011101010 : data_out = 24'b000000110010011110111111;
    16'b0000110011101011 : data_out = 24'b000000110010100010001001;
    16'b0000110011101100 : data_out = 24'b000000110010100101010100;
    16'b0000110011101101 : data_out = 24'b000000110010101000011110;
    16'b0000110011101110 : data_out = 24'b000000110010101011101001;
    16'b0000110011101111 : data_out = 24'b000000110010101110110011;
    16'b0000110011110000 : data_out = 24'b000000110010110001111110;
    16'b0000110011110001 : data_out = 24'b000000110010110101001010;
    16'b0000110011110010 : data_out = 24'b000000110010111000010101;
    16'b0000110011110011 : data_out = 24'b000000110010111011100001;
    16'b0000110011110100 : data_out = 24'b000000110010111110101101;
    16'b0000110011110101 : data_out = 24'b000000110011000001111001;
    16'b0000110011110110 : data_out = 24'b000000110011000101000101;
    16'b0000110011110111 : data_out = 24'b000000110011001000010001;
    16'b0000110011111000 : data_out = 24'b000000110011001011011110;
    16'b0000110011111001 : data_out = 24'b000000110011001110101011;
    16'b0000110011111010 : data_out = 24'b000000110011010001111000;
    16'b0000110011111011 : data_out = 24'b000000110011010101000101;
    16'b0000110011111100 : data_out = 24'b000000110011011000010010;
    16'b0000110011111101 : data_out = 24'b000000110011011011100000;
    16'b0000110011111110 : data_out = 24'b000000110011011110101110;
    16'b0000110011111111 : data_out = 24'b000000110011100001111100;
    16'b0000110100000000 : data_out = 24'b000000110011100101001010;
    16'b0000110100000001 : data_out = 24'b000000110011101000011000;
    16'b0000110100000010 : data_out = 24'b000000110011101011100111;
    16'b0000110100000011 : data_out = 24'b000000110011101110110110;
    16'b0000110100000100 : data_out = 24'b000000110011110010000101;
    16'b0000110100000101 : data_out = 24'b000000110011110101010100;
    16'b0000110100000110 : data_out = 24'b000000110011111000100100;
    16'b0000110100000111 : data_out = 24'b000000110011111011110011;
    16'b0000110100001000 : data_out = 24'b000000110011111111000011;
    16'b0000110100001001 : data_out = 24'b000000110100000010010011;
    16'b0000110100001010 : data_out = 24'b000000110100000101100011;
    16'b0000110100001011 : data_out = 24'b000000110100001000110100;
    16'b0000110100001100 : data_out = 24'b000000110100001100000100;
    16'b0000110100001101 : data_out = 24'b000000110100001111010101;
    16'b0000110100001110 : data_out = 24'b000000110100010010100110;
    16'b0000110100001111 : data_out = 24'b000000110100010101111000;
    16'b0000110100010000 : data_out = 24'b000000110100011001001001;
    16'b0000110100010001 : data_out = 24'b000000110100011100011011;
    16'b0000110100010010 : data_out = 24'b000000110100011111101101;
    16'b0000110100010011 : data_out = 24'b000000110100100010111111;
    16'b0000110100010100 : data_out = 24'b000000110100100110010001;
    16'b0000110100010101 : data_out = 24'b000000110100101001100011;
    16'b0000110100010110 : data_out = 24'b000000110100101100110110;
    16'b0000110100010111 : data_out = 24'b000000110100110000001001;
    16'b0000110100011000 : data_out = 24'b000000110100110011011100;
    16'b0000110100011001 : data_out = 24'b000000110100110110110000;
    16'b0000110100011010 : data_out = 24'b000000110100111010000011;
    16'b0000110100011011 : data_out = 24'b000000110100111101010111;
    16'b0000110100011100 : data_out = 24'b000000110101000000101011;
    16'b0000110100011101 : data_out = 24'b000000110101000011111111;
    16'b0000110100011110 : data_out = 24'b000000110101000111010011;
    16'b0000110100011111 : data_out = 24'b000000110101001010101000;
    16'b0000110100100000 : data_out = 24'b000000110101001101111101;
    16'b0000110100100001 : data_out = 24'b000000110101010001010010;
    16'b0000110100100010 : data_out = 24'b000000110101010100100111;
    16'b0000110100100011 : data_out = 24'b000000110101010111111100;
    16'b0000110100100100 : data_out = 24'b000000110101011011010010;
    16'b0000110100100101 : data_out = 24'b000000110101011110100111;
    16'b0000110100100110 : data_out = 24'b000000110101100001111110;
    16'b0000110100100111 : data_out = 24'b000000110101100101010100;
    16'b0000110100101000 : data_out = 24'b000000110101101000101010;
    16'b0000110100101001 : data_out = 24'b000000110101101100000001;
    16'b0000110100101010 : data_out = 24'b000000110101101111011000;
    16'b0000110100101011 : data_out = 24'b000000110101110010101111;
    16'b0000110100101100 : data_out = 24'b000000110101110110000110;
    16'b0000110100101101 : data_out = 24'b000000110101111001011110;
    16'b0000110100101110 : data_out = 24'b000000110101111100110101;
    16'b0000110100101111 : data_out = 24'b000000110110000000001101;
    16'b0000110100110000 : data_out = 24'b000000110110000011100101;
    16'b0000110100110001 : data_out = 24'b000000110110000110111110;
    16'b0000110100110010 : data_out = 24'b000000110110001010010110;
    16'b0000110100110011 : data_out = 24'b000000110110001101101111;
    16'b0000110100110100 : data_out = 24'b000000110110010001001000;
    16'b0000110100110101 : data_out = 24'b000000110110010100100001;
    16'b0000110100110110 : data_out = 24'b000000110110010111111010;
    16'b0000110100110111 : data_out = 24'b000000110110011011010100;
    16'b0000110100111000 : data_out = 24'b000000110110011110101110;
    16'b0000110100111001 : data_out = 24'b000000110110100010001000;
    16'b0000110100111010 : data_out = 24'b000000110110100101100010;
    16'b0000110100111011 : data_out = 24'b000000110110101000111101;
    16'b0000110100111100 : data_out = 24'b000000110110101100010111;
    16'b0000110100111101 : data_out = 24'b000000110110101111110010;
    16'b0000110100111110 : data_out = 24'b000000110110110011001101;
    16'b0000110100111111 : data_out = 24'b000000110110110110101000;
    16'b0000110101000000 : data_out = 24'b000000110110111010000100;
    16'b0000110101000001 : data_out = 24'b000000110110111101100000;
    16'b0000110101000010 : data_out = 24'b000000110111000000111100;
    16'b0000110101000011 : data_out = 24'b000000110111000100011000;
    16'b0000110101000100 : data_out = 24'b000000110111000111110100;
    16'b0000110101000101 : data_out = 24'b000000110111001011010001;
    16'b0000110101000110 : data_out = 24'b000000110111001110101110;
    16'b0000110101000111 : data_out = 24'b000000110111010010001011;
    16'b0000110101001000 : data_out = 24'b000000110111010101101000;
    16'b0000110101001001 : data_out = 24'b000000110111011001000101;
    16'b0000110101001010 : data_out = 24'b000000110111011100100011;
    16'b0000110101001011 : data_out = 24'b000000110111100000000001;
    16'b0000110101001100 : data_out = 24'b000000110111100011011111;
    16'b0000110101001101 : data_out = 24'b000000110111100110111101;
    16'b0000110101001110 : data_out = 24'b000000110111101010011100;
    16'b0000110101001111 : data_out = 24'b000000110111101101111011;
    16'b0000110101010000 : data_out = 24'b000000110111110001011010;
    16'b0000110101010001 : data_out = 24'b000000110111110100111001;
    16'b0000110101010010 : data_out = 24'b000000110111111000011000;
    16'b0000110101010011 : data_out = 24'b000000110111111011111000;
    16'b0000110101010100 : data_out = 24'b000000110111111111011000;
    16'b0000110101010101 : data_out = 24'b000000111000000010111000;
    16'b0000110101010110 : data_out = 24'b000000111000000110011000;
    16'b0000110101010111 : data_out = 24'b000000111000001001111001;
    16'b0000110101011000 : data_out = 24'b000000111000001101011001;
    16'b0000110101011001 : data_out = 24'b000000111000010000111010;
    16'b0000110101011010 : data_out = 24'b000000111000010100011011;
    16'b0000110101011011 : data_out = 24'b000000111000010111111101;
    16'b0000110101011100 : data_out = 24'b000000111000011011011110;
    16'b0000110101011101 : data_out = 24'b000000111000011111000000;
    16'b0000110101011110 : data_out = 24'b000000111000100010100010;
    16'b0000110101011111 : data_out = 24'b000000111000100110000101;
    16'b0000110101100000 : data_out = 24'b000000111000101001100111;
    16'b0000110101100001 : data_out = 24'b000000111000101101001010;
    16'b0000110101100010 : data_out = 24'b000000111000110000101101;
    16'b0000110101100011 : data_out = 24'b000000111000110100010000;
    16'b0000110101100100 : data_out = 24'b000000111000110111110011;
    16'b0000110101100101 : data_out = 24'b000000111000111011010111;
    16'b0000110101100110 : data_out = 24'b000000111000111110111011;
    16'b0000110101100111 : data_out = 24'b000000111001000010011111;
    16'b0000110101101000 : data_out = 24'b000000111001000110000011;
    16'b0000110101101001 : data_out = 24'b000000111001001001101000;
    16'b0000110101101010 : data_out = 24'b000000111001001101001100;
    16'b0000110101101011 : data_out = 24'b000000111001010000110001;
    16'b0000110101101100 : data_out = 24'b000000111001010100010110;
    16'b0000110101101101 : data_out = 24'b000000111001010111111100;
    16'b0000110101101110 : data_out = 24'b000000111001011011100001;
    16'b0000110101101111 : data_out = 24'b000000111001011111000111;
    16'b0000110101110000 : data_out = 24'b000000111001100010101101;
    16'b0000110101110001 : data_out = 24'b000000111001100110010011;
    16'b0000110101110010 : data_out = 24'b000000111001101001111010;
    16'b0000110101110011 : data_out = 24'b000000111001101101100001;
    16'b0000110101110100 : data_out = 24'b000000111001110001001000;
    16'b0000110101110101 : data_out = 24'b000000111001110100101111;
    16'b0000110101110110 : data_out = 24'b000000111001111000010110;
    16'b0000110101110111 : data_out = 24'b000000111001111011111110;
    16'b0000110101111000 : data_out = 24'b000000111001111111100110;
    16'b0000110101111001 : data_out = 24'b000000111010000011001110;
    16'b0000110101111010 : data_out = 24'b000000111010000110110110;
    16'b0000110101111011 : data_out = 24'b000000111010001010011111;
    16'b0000110101111100 : data_out = 24'b000000111010001110000111;
    16'b0000110101111101 : data_out = 24'b000000111010010001110000;
    16'b0000110101111110 : data_out = 24'b000000111010010101011010;
    16'b0000110101111111 : data_out = 24'b000000111010011001000011;
    16'b0000110110000000 : data_out = 24'b000000111010011100101101;
    16'b0000110110000001 : data_out = 24'b000000111010100000010111;
    16'b0000110110000010 : data_out = 24'b000000111010100100000001;
    16'b0000110110000011 : data_out = 24'b000000111010100111101011;
    16'b0000110110000100 : data_out = 24'b000000111010101011010110;
    16'b0000110110000101 : data_out = 24'b000000111010101111000001;
    16'b0000110110000110 : data_out = 24'b000000111010110010101100;
    16'b0000110110000111 : data_out = 24'b000000111010110110010111;
    16'b0000110110001000 : data_out = 24'b000000111010111010000011;
    16'b0000110110001001 : data_out = 24'b000000111010111101101110;
    16'b0000110110001010 : data_out = 24'b000000111011000001011010;
    16'b0000110110001011 : data_out = 24'b000000111011000101000110;
    16'b0000110110001100 : data_out = 24'b000000111011001000110011;
    16'b0000110110001101 : data_out = 24'b000000111011001100100000;
    16'b0000110110001110 : data_out = 24'b000000111011010000001100;
    16'b0000110110001111 : data_out = 24'b000000111011010011111010;
    16'b0000110110010000 : data_out = 24'b000000111011010111100111;
    16'b0000110110010001 : data_out = 24'b000000111011011011010101;
    16'b0000110110010010 : data_out = 24'b000000111011011111000010;
    16'b0000110110010011 : data_out = 24'b000000111011100010110000;
    16'b0000110110010100 : data_out = 24'b000000111011100110011111;
    16'b0000110110010101 : data_out = 24'b000000111011101010001101;
    16'b0000110110010110 : data_out = 24'b000000111011101101111100;
    16'b0000110110010111 : data_out = 24'b000000111011110001101011;
    16'b0000110110011000 : data_out = 24'b000000111011110101011010;
    16'b0000110110011001 : data_out = 24'b000000111011111001001010;
    16'b0000110110011010 : data_out = 24'b000000111011111100111001;
    16'b0000110110011011 : data_out = 24'b000000111100000000101001;
    16'b0000110110011100 : data_out = 24'b000000111100000100011001;
    16'b0000110110011101 : data_out = 24'b000000111100001000001010;
    16'b0000110110011110 : data_out = 24'b000000111100001011111010;
    16'b0000110110011111 : data_out = 24'b000000111100001111101011;
    16'b0000110110100000 : data_out = 24'b000000111100010011011100;
    16'b0000110110100001 : data_out = 24'b000000111100010111001110;
    16'b0000110110100010 : data_out = 24'b000000111100011010111111;
    16'b0000110110100011 : data_out = 24'b000000111100011110110001;
    16'b0000110110100100 : data_out = 24'b000000111100100010100011;
    16'b0000110110100101 : data_out = 24'b000000111100100110010101;
    16'b0000110110100110 : data_out = 24'b000000111100101010001000;
    16'b0000110110100111 : data_out = 24'b000000111100101101111011;
    16'b0000110110101000 : data_out = 24'b000000111100110001101110;
    16'b0000110110101001 : data_out = 24'b000000111100110101100001;
    16'b0000110110101010 : data_out = 24'b000000111100111001010100;
    16'b0000110110101011 : data_out = 24'b000000111100111101001000;
    16'b0000110110101100 : data_out = 24'b000000111101000000111100;
    16'b0000110110101101 : data_out = 24'b000000111101000100110000;
    16'b0000110110101110 : data_out = 24'b000000111101001000100101;
    16'b0000110110101111 : data_out = 24'b000000111101001100011001;
    16'b0000110110110000 : data_out = 24'b000000111101010000001110;
    16'b0000110110110001 : data_out = 24'b000000111101010100000011;
    16'b0000110110110010 : data_out = 24'b000000111101010111111001;
    16'b0000110110110011 : data_out = 24'b000000111101011011101110;
    16'b0000110110110100 : data_out = 24'b000000111101011111100100;
    16'b0000110110110101 : data_out = 24'b000000111101100011011010;
    16'b0000110110110110 : data_out = 24'b000000111101100111010001;
    16'b0000110110110111 : data_out = 24'b000000111101101011000111;
    16'b0000110110111000 : data_out = 24'b000000111101101110111110;
    16'b0000110110111001 : data_out = 24'b000000111101110010110101;
    16'b0000110110111010 : data_out = 24'b000000111101110110101100;
    16'b0000110110111011 : data_out = 24'b000000111101111010100100;
    16'b0000110110111100 : data_out = 24'b000000111101111110011100;
    16'b0000110110111101 : data_out = 24'b000000111110000010010100;
    16'b0000110110111110 : data_out = 24'b000000111110000110001100;
    16'b0000110110111111 : data_out = 24'b000000111110001010000100;
    16'b0000110111000000 : data_out = 24'b000000111110001101111101;
    16'b0000110111000001 : data_out = 24'b000000111110010001110110;
    16'b0000110111000010 : data_out = 24'b000000111110010101101111;
    16'b0000110111000011 : data_out = 24'b000000111110011001101001;
    16'b0000110111000100 : data_out = 24'b000000111110011101100011;
    16'b0000110111000101 : data_out = 24'b000000111110100001011101;
    16'b0000110111000110 : data_out = 24'b000000111110100101010111;
    16'b0000110111000111 : data_out = 24'b000000111110101001010001;
    16'b0000110111001000 : data_out = 24'b000000111110101101001100;
    16'b0000110111001001 : data_out = 24'b000000111110110001000111;
    16'b0000110111001010 : data_out = 24'b000000111110110101000010;
    16'b0000110111001011 : data_out = 24'b000000111110111000111110;
    16'b0000110111001100 : data_out = 24'b000000111110111100111001;
    16'b0000110111001101 : data_out = 24'b000000111111000000110101;
    16'b0000110111001110 : data_out = 24'b000000111111000100110001;
    16'b0000110111001111 : data_out = 24'b000000111111001000101110;
    16'b0000110111010000 : data_out = 24'b000000111111001100101010;
    16'b0000110111010001 : data_out = 24'b000000111111010000100111;
    16'b0000110111010010 : data_out = 24'b000000111111010100100100;
    16'b0000110111010011 : data_out = 24'b000000111111011000100010;
    16'b0000110111010100 : data_out = 24'b000000111111011100100000;
    16'b0000110111010101 : data_out = 24'b000000111111100000011101;
    16'b0000110111010110 : data_out = 24'b000000111111100100011100;
    16'b0000110111010111 : data_out = 24'b000000111111101000011010;
    16'b0000110111011000 : data_out = 24'b000000111111101100011001;
    16'b0000110111011001 : data_out = 24'b000000111111110000011000;
    16'b0000110111011010 : data_out = 24'b000000111111110100010111;
    16'b0000110111011011 : data_out = 24'b000000111111111000010110;
    16'b0000110111011100 : data_out = 24'b000000111111111100010110;
    16'b0000110111011101 : data_out = 24'b000001000000000000010110;
    16'b0000110111011110 : data_out = 24'b000001000000000100010110;
    16'b0000110111011111 : data_out = 24'b000001000000001000010110;
    16'b0000110111100000 : data_out = 24'b000001000000001100010111;
    16'b0000110111100001 : data_out = 24'b000001000000010000011000;
    16'b0000110111100010 : data_out = 24'b000001000000010100011001;
    16'b0000110111100011 : data_out = 24'b000001000000011000011010;
    16'b0000110111100100 : data_out = 24'b000001000000011100011100;
    16'b0000110111100101 : data_out = 24'b000001000000100000011110;
    16'b0000110111100110 : data_out = 24'b000001000000100100100000;
    16'b0000110111100111 : data_out = 24'b000001000000101000100010;
    16'b0000110111101000 : data_out = 24'b000001000000101100100101;
    16'b0000110111101001 : data_out = 24'b000001000000110000101000;
    16'b0000110111101010 : data_out = 24'b000001000000110100101011;
    16'b0000110111101011 : data_out = 24'b000001000000111000101111;
    16'b0000110111101100 : data_out = 24'b000001000000111100110010;
    16'b0000110111101101 : data_out = 24'b000001000001000000110110;
    16'b0000110111101110 : data_out = 24'b000001000001000100111010;
    16'b0000110111101111 : data_out = 24'b000001000001001000111111;
    16'b0000110111110000 : data_out = 24'b000001000001001101000011;
    16'b0000110111110001 : data_out = 24'b000001000001010001001000;
    16'b0000110111110010 : data_out = 24'b000001000001010101001110;
    16'b0000110111110011 : data_out = 24'b000001000001011001010011;
    16'b0000110111110100 : data_out = 24'b000001000001011101011001;
    16'b0000110111110101 : data_out = 24'b000001000001100001011111;
    16'b0000110111110110 : data_out = 24'b000001000001100101100101;
    16'b0000110111110111 : data_out = 24'b000001000001101001101011;
    16'b0000110111111000 : data_out = 24'b000001000001101101110010;
    16'b0000110111111001 : data_out = 24'b000001000001110001111001;
    16'b0000110111111010 : data_out = 24'b000001000001110110000000;
    16'b0000110111111011 : data_out = 24'b000001000001111010001000;
    16'b0000110111111100 : data_out = 24'b000001000001111110010000;
    16'b0000110111111101 : data_out = 24'b000001000010000010011000;
    16'b0000110111111110 : data_out = 24'b000001000010000110100000;
    16'b0000110111111111 : data_out = 24'b000001000010001010101000;
    16'b0000111000000000 : data_out = 24'b000001000010001110110001;
    16'b0000111000000001 : data_out = 24'b000001000010010010111010;
    16'b0000111000000010 : data_out = 24'b000001000010010111000100;
    16'b0000111000000011 : data_out = 24'b000001000010011011001101;
    16'b0000111000000100 : data_out = 24'b000001000010011111010111;
    16'b0000111000000101 : data_out = 24'b000001000010100011100001;
    16'b0000111000000110 : data_out = 24'b000001000010100111101011;
    16'b0000111000000111 : data_out = 24'b000001000010101011110110;
    16'b0000111000001000 : data_out = 24'b000001000010110000000001;
    16'b0000111000001001 : data_out = 24'b000001000010110100001100;
    16'b0000111000001010 : data_out = 24'b000001000010111000010111;
    16'b0000111000001011 : data_out = 24'b000001000010111100100011;
    16'b0000111000001100 : data_out = 24'b000001000011000000101111;
    16'b0000111000001101 : data_out = 24'b000001000011000100111011;
    16'b0000111000001110 : data_out = 24'b000001000011001001001000;
    16'b0000111000001111 : data_out = 24'b000001000011001101010100;
    16'b0000111000010000 : data_out = 24'b000001000011010001100001;
    16'b0000111000010001 : data_out = 24'b000001000011010101101111;
    16'b0000111000010010 : data_out = 24'b000001000011011001111100;
    16'b0000111000010011 : data_out = 24'b000001000011011110001010;
    16'b0000111000010100 : data_out = 24'b000001000011100010011000;
    16'b0000111000010101 : data_out = 24'b000001000011100110100110;
    16'b0000111000010110 : data_out = 24'b000001000011101010110101;
    16'b0000111000010111 : data_out = 24'b000001000011101111000011;
    16'b0000111000011000 : data_out = 24'b000001000011110011010011;
    16'b0000111000011001 : data_out = 24'b000001000011110111100010;
    16'b0000111000011010 : data_out = 24'b000001000011111011110001;
    16'b0000111000011011 : data_out = 24'b000001000100000000000001;
    16'b0000111000011100 : data_out = 24'b000001000100000100010001;
    16'b0000111000011101 : data_out = 24'b000001000100001000100010;
    16'b0000111000011110 : data_out = 24'b000001000100001100110011;
    16'b0000111000011111 : data_out = 24'b000001000100010001000011;
    16'b0000111000100000 : data_out = 24'b000001000100010101010101;
    16'b0000111000100001 : data_out = 24'b000001000100011001100110;
    16'b0000111000100010 : data_out = 24'b000001000100011101111000;
    16'b0000111000100011 : data_out = 24'b000001000100100010001010;
    16'b0000111000100100 : data_out = 24'b000001000100100110011100;
    16'b0000111000100101 : data_out = 24'b000001000100101010101111;
    16'b0000111000100110 : data_out = 24'b000001000100101111000010;
    16'b0000111000100111 : data_out = 24'b000001000100110011010101;
    16'b0000111000101000 : data_out = 24'b000001000100110111101000;
    16'b0000111000101001 : data_out = 24'b000001000100111011111100;
    16'b0000111000101010 : data_out = 24'b000001000101000000001111;
    16'b0000111000101011 : data_out = 24'b000001000101000100100100;
    16'b0000111000101100 : data_out = 24'b000001000101001000111000;
    16'b0000111000101101 : data_out = 24'b000001000101001101001101;
    16'b0000111000101110 : data_out = 24'b000001000101010001100010;
    16'b0000111000101111 : data_out = 24'b000001000101010101110111;
    16'b0000111000110000 : data_out = 24'b000001000101011010001100;
    16'b0000111000110001 : data_out = 24'b000001000101011110100010;
    16'b0000111000110010 : data_out = 24'b000001000101100010111000;
    16'b0000111000110011 : data_out = 24'b000001000101100111001111;
    16'b0000111000110100 : data_out = 24'b000001000101101011100101;
    16'b0000111000110101 : data_out = 24'b000001000101101111111100;
    16'b0000111000110110 : data_out = 24'b000001000101110100010011;
    16'b0000111000110111 : data_out = 24'b000001000101111000101010;
    16'b0000111000111000 : data_out = 24'b000001000101111101000010;
    16'b0000111000111001 : data_out = 24'b000001000110000001011010;
    16'b0000111000111010 : data_out = 24'b000001000110000101110010;
    16'b0000111000111011 : data_out = 24'b000001000110001010001011;
    16'b0000111000111100 : data_out = 24'b000001000110001110100100;
    16'b0000111000111101 : data_out = 24'b000001000110010010111101;
    16'b0000111000111110 : data_out = 24'b000001000110010111010110;
    16'b0000111000111111 : data_out = 24'b000001000110011011110000;
    16'b0000111001000000 : data_out = 24'b000001000110100000001001;
    16'b0000111001000001 : data_out = 24'b000001000110100100100100;
    16'b0000111001000010 : data_out = 24'b000001000110101000111110;
    16'b0000111001000011 : data_out = 24'b000001000110101101011001;
    16'b0000111001000100 : data_out = 24'b000001000110110001110100;
    16'b0000111001000101 : data_out = 24'b000001000110110110001111;
    16'b0000111001000110 : data_out = 24'b000001000110111010101010;
    16'b0000111001000111 : data_out = 24'b000001000110111111000110;
    16'b0000111001001000 : data_out = 24'b000001000111000011100010;
    16'b0000111001001001 : data_out = 24'b000001000111000111111111;
    16'b0000111001001010 : data_out = 24'b000001000111001100011011;
    16'b0000111001001011 : data_out = 24'b000001000111010000111000;
    16'b0000111001001100 : data_out = 24'b000001000111010101010101;
    16'b0000111001001101 : data_out = 24'b000001000111011001110011;
    16'b0000111001001110 : data_out = 24'b000001000111011110010001;
    16'b0000111001001111 : data_out = 24'b000001000111100010101111;
    16'b0000111001010000 : data_out = 24'b000001000111100111001101;
    16'b0000111001010001 : data_out = 24'b000001000111101011101100;
    16'b0000111001010010 : data_out = 24'b000001000111110000001011;
    16'b0000111001010011 : data_out = 24'b000001000111110100101010;
    16'b0000111001010100 : data_out = 24'b000001000111111001001001;
    16'b0000111001010101 : data_out = 24'b000001000111111101101001;
    16'b0000111001010110 : data_out = 24'b000001001000000010001001;
    16'b0000111001010111 : data_out = 24'b000001001000000110101001;
    16'b0000111001011000 : data_out = 24'b000001001000001011001010;
    16'b0000111001011001 : data_out = 24'b000001001000001111101010;
    16'b0000111001011010 : data_out = 24'b000001001000010100001100;
    16'b0000111001011011 : data_out = 24'b000001001000011000101101;
    16'b0000111001011100 : data_out = 24'b000001001000011101001111;
    16'b0000111001011101 : data_out = 24'b000001001000100001110001;
    16'b0000111001011110 : data_out = 24'b000001001000100110010011;
    16'b0000111001011111 : data_out = 24'b000001001000101010110101;
    16'b0000111001100000 : data_out = 24'b000001001000101111011000;
    16'b0000111001100001 : data_out = 24'b000001001000110011111011;
    16'b0000111001100010 : data_out = 24'b000001001000111000011111;
    16'b0000111001100011 : data_out = 24'b000001001000111101000010;
    16'b0000111001100100 : data_out = 24'b000001001001000001100110;
    16'b0000111001100101 : data_out = 24'b000001001001000110001011;
    16'b0000111001100110 : data_out = 24'b000001001001001010101111;
    16'b0000111001100111 : data_out = 24'b000001001001001111010100;
    16'b0000111001101000 : data_out = 24'b000001001001010011111001;
    16'b0000111001101001 : data_out = 24'b000001001001011000011110;
    16'b0000111001101010 : data_out = 24'b000001001001011101000100;
    16'b0000111001101011 : data_out = 24'b000001001001100001101010;
    16'b0000111001101100 : data_out = 24'b000001001001100110010000;
    16'b0000111001101101 : data_out = 24'b000001001001101010110111;
    16'b0000111001101110 : data_out = 24'b000001001001101111011110;
    16'b0000111001101111 : data_out = 24'b000001001001110100000101;
    16'b0000111001110000 : data_out = 24'b000001001001111000101100;
    16'b0000111001110001 : data_out = 24'b000001001001111101010100;
    16'b0000111001110010 : data_out = 24'b000001001010000001111100;
    16'b0000111001110011 : data_out = 24'b000001001010000110100100;
    16'b0000111001110100 : data_out = 24'b000001001010001011001101;
    16'b0000111001110101 : data_out = 24'b000001001010001111110110;
    16'b0000111001110110 : data_out = 24'b000001001010010100011111;
    16'b0000111001110111 : data_out = 24'b000001001010011001001000;
    16'b0000111001111000 : data_out = 24'b000001001010011101110010;
    16'b0000111001111001 : data_out = 24'b000001001010100010011100;
    16'b0000111001111010 : data_out = 24'b000001001010100111000110;
    16'b0000111001111011 : data_out = 24'b000001001010101011110001;
    16'b0000111001111100 : data_out = 24'b000001001010110000011100;
    16'b0000111001111101 : data_out = 24'b000001001010110101000111;
    16'b0000111001111110 : data_out = 24'b000001001010111001110010;
    16'b0000111001111111 : data_out = 24'b000001001010111110011110;
    16'b0000111010000000 : data_out = 24'b000001001011000011001010;
    16'b0000111010000001 : data_out = 24'b000001001011000111110110;
    16'b0000111010000010 : data_out = 24'b000001001011001100100011;
    16'b0000111010000011 : data_out = 24'b000001001011010001010000;
    16'b0000111010000100 : data_out = 24'b000001001011010101111101;
    16'b0000111010000101 : data_out = 24'b000001001011011010101011;
    16'b0000111010000110 : data_out = 24'b000001001011011111011001;
    16'b0000111010000111 : data_out = 24'b000001001011100100000111;
    16'b0000111010001000 : data_out = 24'b000001001011101000110101;
    16'b0000111010001001 : data_out = 24'b000001001011101101100100;
    16'b0000111010001010 : data_out = 24'b000001001011110010010011;
    16'b0000111010001011 : data_out = 24'b000001001011110111000010;
    16'b0000111010001100 : data_out = 24'b000001001011111011110010;
    16'b0000111010001101 : data_out = 24'b000001001100000000100001;
    16'b0000111010001110 : data_out = 24'b000001001100000101010010;
    16'b0000111010001111 : data_out = 24'b000001001100001010000010;
    16'b0000111010010000 : data_out = 24'b000001001100001110110011;
    16'b0000111010010001 : data_out = 24'b000001001100010011100100;
    16'b0000111010010010 : data_out = 24'b000001001100011000010101;
    16'b0000111010010011 : data_out = 24'b000001001100011101000111;
    16'b0000111010010100 : data_out = 24'b000001001100100001111001;
    16'b0000111010010101 : data_out = 24'b000001001100100110101011;
    16'b0000111010010110 : data_out = 24'b000001001100101011011110;
    16'b0000111010010111 : data_out = 24'b000001001100110000010001;
    16'b0000111010011000 : data_out = 24'b000001001100110101000100;
    16'b0000111010011001 : data_out = 24'b000001001100111001110111;
    16'b0000111010011010 : data_out = 24'b000001001100111110101011;
    16'b0000111010011011 : data_out = 24'b000001001101000011011111;
    16'b0000111010011100 : data_out = 24'b000001001101001000010100;
    16'b0000111010011101 : data_out = 24'b000001001101001101001000;
    16'b0000111010011110 : data_out = 24'b000001001101010001111101;
    16'b0000111010011111 : data_out = 24'b000001001101010110110010;
    16'b0000111010100000 : data_out = 24'b000001001101011011101000;
    16'b0000111010100001 : data_out = 24'b000001001101100000011110;
    16'b0000111010100010 : data_out = 24'b000001001101100101010100;
    16'b0000111010100011 : data_out = 24'b000001001101101010001011;
    16'b0000111010100100 : data_out = 24'b000001001101101111000001;
    16'b0000111010100101 : data_out = 24'b000001001101110011111000;
    16'b0000111010100110 : data_out = 24'b000001001101111000110000;
    16'b0000111010100111 : data_out = 24'b000001001101111101101000;
    16'b0000111010101000 : data_out = 24'b000001001110000010100000;
    16'b0000111010101001 : data_out = 24'b000001001110000111011000;
    16'b0000111010101010 : data_out = 24'b000001001110001100010000;
    16'b0000111010101011 : data_out = 24'b000001001110010001001001;
    16'b0000111010101100 : data_out = 24'b000001001110010110000011;
    16'b0000111010101101 : data_out = 24'b000001001110011010111100;
    16'b0000111010101110 : data_out = 24'b000001001110011111110110;
    16'b0000111010101111 : data_out = 24'b000001001110100100110000;
    16'b0000111010110000 : data_out = 24'b000001001110101001101011;
    16'b0000111010110001 : data_out = 24'b000001001110101110100101;
    16'b0000111010110010 : data_out = 24'b000001001110110011100000;
    16'b0000111010110011 : data_out = 24'b000001001110111000011100;
    16'b0000111010110100 : data_out = 24'b000001001110111101010111;
    16'b0000111010110101 : data_out = 24'b000001001111000010010011;
    16'b0000111010110110 : data_out = 24'b000001001111000111010000;
    16'b0000111010110111 : data_out = 24'b000001001111001100001100;
    16'b0000111010111000 : data_out = 24'b000001001111010001001001;
    16'b0000111010111001 : data_out = 24'b000001001111010110000111;
    16'b0000111010111010 : data_out = 24'b000001001111011011000100;
    16'b0000111010111011 : data_out = 24'b000001001111100000000010;
    16'b0000111010111100 : data_out = 24'b000001001111100101000000;
    16'b0000111010111101 : data_out = 24'b000001001111101001111111;
    16'b0000111010111110 : data_out = 24'b000001001111101110111101;
    16'b0000111010111111 : data_out = 24'b000001001111110011111100;
    16'b0000111011000000 : data_out = 24'b000001001111111000111100;
    16'b0000111011000001 : data_out = 24'b000001001111111101111100;
    16'b0000111011000010 : data_out = 24'b000001010000000010111100;
    16'b0000111011000011 : data_out = 24'b000001010000000111111100;
    16'b0000111011000100 : data_out = 24'b000001010000001100111101;
    16'b0000111011000101 : data_out = 24'b000001010000010001111101;
    16'b0000111011000110 : data_out = 24'b000001010000010110111111;
    16'b0000111011000111 : data_out = 24'b000001010000011100000000;
    16'b0000111011001000 : data_out = 24'b000001010000100001000010;
    16'b0000111011001001 : data_out = 24'b000001010000100110000100;
    16'b0000111011001010 : data_out = 24'b000001010000101011000111;
    16'b0000111011001011 : data_out = 24'b000001010000110000001010;
    16'b0000111011001100 : data_out = 24'b000001010000110101001101;
    16'b0000111011001101 : data_out = 24'b000001010000111010010001;
    16'b0000111011001110 : data_out = 24'b000001010000111111010100;
    16'b0000111011001111 : data_out = 24'b000001010001000100011000;
    16'b0000111011010000 : data_out = 24'b000001010001001001011101;
    16'b0000111011010001 : data_out = 24'b000001010001001110100010;
    16'b0000111011010010 : data_out = 24'b000001010001010011100111;
    16'b0000111011010011 : data_out = 24'b000001010001011000101100;
    16'b0000111011010100 : data_out = 24'b000001010001011101110010;
    16'b0000111011010101 : data_out = 24'b000001010001100010111000;
    16'b0000111011010110 : data_out = 24'b000001010001100111111110;
    16'b0000111011010111 : data_out = 24'b000001010001101101000101;
    16'b0000111011011000 : data_out = 24'b000001010001110010001100;
    16'b0000111011011001 : data_out = 24'b000001010001110111010011;
    16'b0000111011011010 : data_out = 24'b000001010001111100011011;
    16'b0000111011011011 : data_out = 24'b000001010010000001100011;
    16'b0000111011011100 : data_out = 24'b000001010010000110101011;
    16'b0000111011011101 : data_out = 24'b000001010010001011110011;
    16'b0000111011011110 : data_out = 24'b000001010010010000111100;
    16'b0000111011011111 : data_out = 24'b000001010010010110000110;
    16'b0000111011100000 : data_out = 24'b000001010010011011001111;
    16'b0000111011100001 : data_out = 24'b000001010010100000011001;
    16'b0000111011100010 : data_out = 24'b000001010010100101100011;
    16'b0000111011100011 : data_out = 24'b000001010010101010101110;
    16'b0000111011100100 : data_out = 24'b000001010010101111111001;
    16'b0000111011100101 : data_out = 24'b000001010010110101000100;
    16'b0000111011100110 : data_out = 24'b000001010010111010001111;
    16'b0000111011100111 : data_out = 24'b000001010010111111011011;
    16'b0000111011101000 : data_out = 24'b000001010011000100100111;
    16'b0000111011101001 : data_out = 24'b000001010011001001110100;
    16'b0000111011101010 : data_out = 24'b000001010011001111000000;
    16'b0000111011101011 : data_out = 24'b000001010011010100001101;
    16'b0000111011101100 : data_out = 24'b000001010011011001011011;
    16'b0000111011101101 : data_out = 24'b000001010011011110101001;
    16'b0000111011101110 : data_out = 24'b000001010011100011110111;
    16'b0000111011101111 : data_out = 24'b000001010011101001000101;
    16'b0000111011110000 : data_out = 24'b000001010011101110010100;
    16'b0000111011110001 : data_out = 24'b000001010011110011100011;
    16'b0000111011110010 : data_out = 24'b000001010011111000110010;
    16'b0000111011110011 : data_out = 24'b000001010011111110000010;
    16'b0000111011110100 : data_out = 24'b000001010100000011010010;
    16'b0000111011110101 : data_out = 24'b000001010100001000100010;
    16'b0000111011110110 : data_out = 24'b000001010100001101110011;
    16'b0000111011110111 : data_out = 24'b000001010100010011000100;
    16'b0000111011111000 : data_out = 24'b000001010100011000010101;
    16'b0000111011111001 : data_out = 24'b000001010100011101100111;
    16'b0000111011111010 : data_out = 24'b000001010100100010111001;
    16'b0000111011111011 : data_out = 24'b000001010100101000001100;
    16'b0000111011111100 : data_out = 24'b000001010100101101011110;
    16'b0000111011111101 : data_out = 24'b000001010100110010110001;
    16'b0000111011111110 : data_out = 24'b000001010100111000000101;
    16'b0000111011111111 : data_out = 24'b000001010100111101011000;
    16'b0000111100000000 : data_out = 24'b000001010101000010101100;
    16'b0000111100000001 : data_out = 24'b000001010101001000000001;
    16'b0000111100000010 : data_out = 24'b000001010101001101010101;
    16'b0000111100000011 : data_out = 24'b000001010101010010101010;
    16'b0000111100000100 : data_out = 24'b000001010101011000000000;
    16'b0000111100000101 : data_out = 24'b000001010101011101010101;
    16'b0000111100000110 : data_out = 24'b000001010101100010101011;
    16'b0000111100000111 : data_out = 24'b000001010101101000000010;
    16'b0000111100001000 : data_out = 24'b000001010101101101011000;
    16'b0000111100001001 : data_out = 24'b000001010101110010101111;
    16'b0000111100001010 : data_out = 24'b000001010101111000000111;
    16'b0000111100001011 : data_out = 24'b000001010101111101011110;
    16'b0000111100001100 : data_out = 24'b000001010110000010110110;
    16'b0000111100001101 : data_out = 24'b000001010110001000001111;
    16'b0000111100001110 : data_out = 24'b000001010110001101100111;
    16'b0000111100001111 : data_out = 24'b000001010110010011000000;
    16'b0000111100010000 : data_out = 24'b000001010110011000011010;
    16'b0000111100010001 : data_out = 24'b000001010110011101110011;
    16'b0000111100010010 : data_out = 24'b000001010110100011001101;
    16'b0000111100010011 : data_out = 24'b000001010110101000101000;
    16'b0000111100010100 : data_out = 24'b000001010110101110000010;
    16'b0000111100010101 : data_out = 24'b000001010110110011011101;
    16'b0000111100010110 : data_out = 24'b000001010110111000111001;
    16'b0000111100010111 : data_out = 24'b000001010110111110010101;
    16'b0000111100011000 : data_out = 24'b000001010111000011110001;
    16'b0000111100011001 : data_out = 24'b000001010111001001001101;
    16'b0000111100011010 : data_out = 24'b000001010111001110101010;
    16'b0000111100011011 : data_out = 24'b000001010111010100000111;
    16'b0000111100011100 : data_out = 24'b000001010111011001100100;
    16'b0000111100011101 : data_out = 24'b000001010111011111000010;
    16'b0000111100011110 : data_out = 24'b000001010111100100100000;
    16'b0000111100011111 : data_out = 24'b000001010111101001111111;
    16'b0000111100100000 : data_out = 24'b000001010111101111011101;
    16'b0000111100100001 : data_out = 24'b000001010111110100111101;
    16'b0000111100100010 : data_out = 24'b000001010111111010011100;
    16'b0000111100100011 : data_out = 24'b000001010111111111111100;
    16'b0000111100100100 : data_out = 24'b000001011000000101011100;
    16'b0000111100100101 : data_out = 24'b000001011000001010111101;
    16'b0000111100100110 : data_out = 24'b000001011000010000011101;
    16'b0000111100100111 : data_out = 24'b000001011000010101111111;
    16'b0000111100101000 : data_out = 24'b000001011000011011100000;
    16'b0000111100101001 : data_out = 24'b000001011000100001000010;
    16'b0000111100101010 : data_out = 24'b000001011000100110100100;
    16'b0000111100101011 : data_out = 24'b000001011000101100000111;
    16'b0000111100101100 : data_out = 24'b000001011000110001101010;
    16'b0000111100101101 : data_out = 24'b000001011000110111001101;
    16'b0000111100101110 : data_out = 24'b000001011000111100110001;
    16'b0000111100101111 : data_out = 24'b000001011001000010010101;
    16'b0000111100110000 : data_out = 24'b000001011001000111111001;
    16'b0000111100110001 : data_out = 24'b000001011001001101011110;
    16'b0000111100110010 : data_out = 24'b000001011001010011000011;
    16'b0000111100110011 : data_out = 24'b000001011001011000101000;
    16'b0000111100110100 : data_out = 24'b000001011001011110001110;
    16'b0000111100110101 : data_out = 24'b000001011001100011110100;
    16'b0000111100110110 : data_out = 24'b000001011001101001011010;
    16'b0000111100110111 : data_out = 24'b000001011001101111000001;
    16'b0000111100111000 : data_out = 24'b000001011001110100101000;
    16'b0000111100111001 : data_out = 24'b000001011001111010010000;
    16'b0000111100111010 : data_out = 24'b000001011001111111110111;
    16'b0000111100111011 : data_out = 24'b000001011010000101100000;
    16'b0000111100111100 : data_out = 24'b000001011010001011001000;
    16'b0000111100111101 : data_out = 24'b000001011010010000110001;
    16'b0000111100111110 : data_out = 24'b000001011010010110011010;
    16'b0000111100111111 : data_out = 24'b000001011010011100000100;
    16'b0000111101000000 : data_out = 24'b000001011010100001101110;
    16'b0000111101000001 : data_out = 24'b000001011010100111011000;
    16'b0000111101000010 : data_out = 24'b000001011010101101000011;
    16'b0000111101000011 : data_out = 24'b000001011010110010101110;
    16'b0000111101000100 : data_out = 24'b000001011010111000011001;
    16'b0000111101000101 : data_out = 24'b000001011010111110000101;
    16'b0000111101000110 : data_out = 24'b000001011011000011110001;
    16'b0000111101000111 : data_out = 24'b000001011011001001011101;
    16'b0000111101001000 : data_out = 24'b000001011011001111001010;
    16'b0000111101001001 : data_out = 24'b000001011011010100110111;
    16'b0000111101001010 : data_out = 24'b000001011011011010100101;
    16'b0000111101001011 : data_out = 24'b000001011011100000010010;
    16'b0000111101001100 : data_out = 24'b000001011011100110000001;
    16'b0000111101001101 : data_out = 24'b000001011011101011101111;
    16'b0000111101001110 : data_out = 24'b000001011011110001011110;
    16'b0000111101001111 : data_out = 24'b000001011011110111001101;
    16'b0000111101010000 : data_out = 24'b000001011011111100111101;
    16'b0000111101010001 : data_out = 24'b000001011100000010101101;
    16'b0000111101010010 : data_out = 24'b000001011100001000011101;
    16'b0000111101010011 : data_out = 24'b000001011100001110001110;
    16'b0000111101010100 : data_out = 24'b000001011100010011111111;
    16'b0000111101010101 : data_out = 24'b000001011100011001110001;
    16'b0000111101010110 : data_out = 24'b000001011100011111100010;
    16'b0000111101010111 : data_out = 24'b000001011100100101010100;
    16'b0000111101011000 : data_out = 24'b000001011100101011000111;
    16'b0000111101011001 : data_out = 24'b000001011100110000111010;
    16'b0000111101011010 : data_out = 24'b000001011100110110101101;
    16'b0000111101011011 : data_out = 24'b000001011100111100100001;
    16'b0000111101011100 : data_out = 24'b000001011101000010010101;
    16'b0000111101011101 : data_out = 24'b000001011101001000001001;
    16'b0000111101011110 : data_out = 24'b000001011101001101111110;
    16'b0000111101011111 : data_out = 24'b000001011101010011110011;
    16'b0000111101100000 : data_out = 24'b000001011101011001101000;
    16'b0000111101100001 : data_out = 24'b000001011101011111011110;
    16'b0000111101100010 : data_out = 24'b000001011101100101010100;
    16'b0000111101100011 : data_out = 24'b000001011101101011001011;
    16'b0000111101100100 : data_out = 24'b000001011101110001000001;
    16'b0000111101100101 : data_out = 24'b000001011101110110111001;
    16'b0000111101100110 : data_out = 24'b000001011101111100110000;
    16'b0000111101100111 : data_out = 24'b000001011110000010101000;
    16'b0000111101101000 : data_out = 24'b000001011110001000100001;
    16'b0000111101101001 : data_out = 24'b000001011110001110011001;
    16'b0000111101101010 : data_out = 24'b000001011110010100010010;
    16'b0000111101101011 : data_out = 24'b000001011110011010001100;
    16'b0000111101101100 : data_out = 24'b000001011110100000000110;
    16'b0000111101101101 : data_out = 24'b000001011110100110000000;
    16'b0000111101101110 : data_out = 24'b000001011110101011111010;
    16'b0000111101101111 : data_out = 24'b000001011110110001110101;
    16'b0000111101110000 : data_out = 24'b000001011110110111110001;
    16'b0000111101110001 : data_out = 24'b000001011110111101101100;
    16'b0000111101110010 : data_out = 24'b000001011111000011101000;
    16'b0000111101110011 : data_out = 24'b000001011111001001100101;
    16'b0000111101110100 : data_out = 24'b000001011111001111100010;
    16'b0000111101110101 : data_out = 24'b000001011111010101011111;
    16'b0000111101110110 : data_out = 24'b000001011111011011011100;
    16'b0000111101110111 : data_out = 24'b000001011111100001011010;
    16'b0000111101111000 : data_out = 24'b000001011111100111011000;
    16'b0000111101111001 : data_out = 24'b000001011111101101010111;
    16'b0000111101111010 : data_out = 24'b000001011111110011010110;
    16'b0000111101111011 : data_out = 24'b000001011111111001010110;
    16'b0000111101111100 : data_out = 24'b000001011111111111010101;
    16'b0000111101111101 : data_out = 24'b000001100000000101010101;
    16'b0000111101111110 : data_out = 24'b000001100000001011010110;
    16'b0000111101111111 : data_out = 24'b000001100000010001010111;
    16'b0000111110000000 : data_out = 24'b000001100000010111011000;
    16'b0000111110000001 : data_out = 24'b000001100000011101011010;
    16'b0000111110000010 : data_out = 24'b000001100000100011011100;
    16'b0000111110000011 : data_out = 24'b000001100000101001011110;
    16'b0000111110000100 : data_out = 24'b000001100000101111100001;
    16'b0000111110000101 : data_out = 24'b000001100000110101100100;
    16'b0000111110000110 : data_out = 24'b000001100000111011101000;
    16'b0000111110000111 : data_out = 24'b000001100001000001101100;
    16'b0000111110001000 : data_out = 24'b000001100001000111110000;
    16'b0000111110001001 : data_out = 24'b000001100001001101110101;
    16'b0000111110001010 : data_out = 24'b000001100001010011111010;
    16'b0000111110001011 : data_out = 24'b000001100001011001111111;
    16'b0000111110001100 : data_out = 24'b000001100001100000000101;
    16'b0000111110001101 : data_out = 24'b000001100001100110001011;
    16'b0000111110001110 : data_out = 24'b000001100001101100010010;
    16'b0000111110001111 : data_out = 24'b000001100001110010011001;
    16'b0000111110010000 : data_out = 24'b000001100001111000100000;
    16'b0000111110010001 : data_out = 24'b000001100001111110101000;
    16'b0000111110010010 : data_out = 24'b000001100010000100110000;
    16'b0000111110010011 : data_out = 24'b000001100010001010111000;
    16'b0000111110010100 : data_out = 24'b000001100010010001000001;
    16'b0000111110010101 : data_out = 24'b000001100010010111001010;
    16'b0000111110010110 : data_out = 24'b000001100010011101010100;
    16'b0000111110010111 : data_out = 24'b000001100010100011011110;
    16'b0000111110011000 : data_out = 24'b000001100010101001101001;
    16'b0000111110011001 : data_out = 24'b000001100010101111110011;
    16'b0000111110011010 : data_out = 24'b000001100010110101111110;
    16'b0000111110011011 : data_out = 24'b000001100010111100001010;
    16'b0000111110011100 : data_out = 24'b000001100011000010010110;
    16'b0000111110011101 : data_out = 24'b000001100011001000100010;
    16'b0000111110011110 : data_out = 24'b000001100011001110101111;
    16'b0000111110011111 : data_out = 24'b000001100011010100111100;
    16'b0000111110100000 : data_out = 24'b000001100011011011001010;
    16'b0000111110100001 : data_out = 24'b000001100011100001011000;
    16'b0000111110100010 : data_out = 24'b000001100011100111100110;
    16'b0000111110100011 : data_out = 24'b000001100011101101110101;
    16'b0000111110100100 : data_out = 24'b000001100011110100000100;
    16'b0000111110100101 : data_out = 24'b000001100011111010010011;
    16'b0000111110100110 : data_out = 24'b000001100100000000100011;
    16'b0000111110100111 : data_out = 24'b000001100100000110110011;
    16'b0000111110101000 : data_out = 24'b000001100100001101000100;
    16'b0000111110101001 : data_out = 24'b000001100100010011010101;
    16'b0000111110101010 : data_out = 24'b000001100100011001100110;
    16'b0000111110101011 : data_out = 24'b000001100100011111111000;
    16'b0000111110101100 : data_out = 24'b000001100100100110001010;
    16'b0000111110101101 : data_out = 24'b000001100100101100011101;
    16'b0000111110101110 : data_out = 24'b000001100100110010110000;
    16'b0000111110101111 : data_out = 24'b000001100100111001000011;
    16'b0000111110110000 : data_out = 24'b000001100100111111010111;
    16'b0000111110110001 : data_out = 24'b000001100101000101101011;
    16'b0000111110110010 : data_out = 24'b000001100101001100000000;
    16'b0000111110110011 : data_out = 24'b000001100101010010010100;
    16'b0000111110110100 : data_out = 24'b000001100101011000101010;
    16'b0000111110110101 : data_out = 24'b000001100101011111000000;
    16'b0000111110110110 : data_out = 24'b000001100101100101010110;
    16'b0000111110110111 : data_out = 24'b000001100101101011101100;
    16'b0000111110111000 : data_out = 24'b000001100101110010000011;
    16'b0000111110111001 : data_out = 24'b000001100101111000011010;
    16'b0000111110111010 : data_out = 24'b000001100101111110110010;
    16'b0000111110111011 : data_out = 24'b000001100110000101001010;
    16'b0000111110111100 : data_out = 24'b000001100110001011100011;
    16'b0000111110111101 : data_out = 24'b000001100110010001111100;
    16'b0000111110111110 : data_out = 24'b000001100110011000010101;
    16'b0000111110111111 : data_out = 24'b000001100110011110101111;
    16'b0000111111000000 : data_out = 24'b000001100110100101001001;
    16'b0000111111000001 : data_out = 24'b000001100110101011100011;
    16'b0000111111000010 : data_out = 24'b000001100110110001111110;
    16'b0000111111000011 : data_out = 24'b000001100110111000011010;
    16'b0000111111000100 : data_out = 24'b000001100110111110110101;
    16'b0000111111000101 : data_out = 24'b000001100111000101010010;
    16'b0000111111000110 : data_out = 24'b000001100111001011101110;
    16'b0000111111000111 : data_out = 24'b000001100111010010001011;
    16'b0000111111001000 : data_out = 24'b000001100111011000101000;
    16'b0000111111001001 : data_out = 24'b000001100111011111000110;
    16'b0000111111001010 : data_out = 24'b000001100111100101100100;
    16'b0000111111001011 : data_out = 24'b000001100111101100000011;
    16'b0000111111001100 : data_out = 24'b000001100111110010100010;
    16'b0000111111001101 : data_out = 24'b000001100111111001000001;
    16'b0000111111001110 : data_out = 24'b000001100111111111100001;
    16'b0000111111001111 : data_out = 24'b000001101000000110000001;
    16'b0000111111010000 : data_out = 24'b000001101000001100100010;
    16'b0000111111010001 : data_out = 24'b000001101000010011000011;
    16'b0000111111010010 : data_out = 24'b000001101000011001100100;
    16'b0000111111010011 : data_out = 24'b000001101000100000000110;
    16'b0000111111010100 : data_out = 24'b000001101000100110101000;
    16'b0000111111010101 : data_out = 24'b000001101000101101001011;
    16'b0000111111010110 : data_out = 24'b000001101000110011101110;
    16'b0000111111010111 : data_out = 24'b000001101000111010010001;
    16'b0000111111011000 : data_out = 24'b000001101001000000110101;
    16'b0000111111011001 : data_out = 24'b000001101001000111011001;
    16'b0000111111011010 : data_out = 24'b000001101001001101111110;
    16'b0000111111011011 : data_out = 24'b000001101001010100100011;
    16'b0000111111011100 : data_out = 24'b000001101001011011001000;
    16'b0000111111011101 : data_out = 24'b000001101001100001101110;
    16'b0000111111011110 : data_out = 24'b000001101001101000010101;
    16'b0000111111011111 : data_out = 24'b000001101001101110111011;
    16'b0000111111100000 : data_out = 24'b000001101001110101100011;
    16'b0000111111100001 : data_out = 24'b000001101001111100001010;
    16'b0000111111100010 : data_out = 24'b000001101010000010110010;
    16'b0000111111100011 : data_out = 24'b000001101010001001011010;
    16'b0000111111100100 : data_out = 24'b000001101010010000000011;
    16'b0000111111100101 : data_out = 24'b000001101010010110101100;
    16'b0000111111100110 : data_out = 24'b000001101010011101010110;
    16'b0000111111100111 : data_out = 24'b000001101010100100000000;
    16'b0000111111101000 : data_out = 24'b000001101010101010101011;
    16'b0000111111101001 : data_out = 24'b000001101010110001010101;
    16'b0000111111101010 : data_out = 24'b000001101010111000000001;
    16'b0000111111101011 : data_out = 24'b000001101010111110101100;
    16'b0000111111101100 : data_out = 24'b000001101011000101011001;
    16'b0000111111101101 : data_out = 24'b000001101011001100000101;
    16'b0000111111101110 : data_out = 24'b000001101011010010110010;
    16'b0000111111101111 : data_out = 24'b000001101011011001011111;
    16'b0000111111110000 : data_out = 24'b000001101011100000001101;
    16'b0000111111110001 : data_out = 24'b000001101011100110111100;
    16'b0000111111110010 : data_out = 24'b000001101011101101101010;
    16'b0000111111110011 : data_out = 24'b000001101011110100011001;
    16'b0000111111110100 : data_out = 24'b000001101011111011001001;
    16'b0000111111110101 : data_out = 24'b000001101100000001111001;
    16'b0000111111110110 : data_out = 24'b000001101100001000101001;
    16'b0000111111110111 : data_out = 24'b000001101100001111011010;
    16'b0000111111111000 : data_out = 24'b000001101100010110001011;
    16'b0000111111111001 : data_out = 24'b000001101100011100111100;
    16'b0000111111111010 : data_out = 24'b000001101100100011101110;
    16'b0000111111111011 : data_out = 24'b000001101100101010100001;
    16'b0000111111111100 : data_out = 24'b000001101100110001010100;
    16'b0000111111111101 : data_out = 24'b000001101100111000000111;
    16'b0000111111111110 : data_out = 24'b000001101100111110111011;
    16'b0000111111111111 : data_out = 24'b000001101101000101101111;
    16'b0001000000000000 : data_out = 24'b000001101101001100100100;
    16'b0001000000000001 : data_out = 24'b000001101101010011011001;
    16'b0001000000000010 : data_out = 24'b000001101101011010001110;
    16'b0001000000000011 : data_out = 24'b000001101101100001000100;
    16'b0001000000000100 : data_out = 24'b000001101101100111111010;
    16'b0001000000000101 : data_out = 24'b000001101101101110110001;
    16'b0001000000000110 : data_out = 24'b000001101101110101101000;
    16'b0001000000000111 : data_out = 24'b000001101101111100100000;
    16'b0001000000001000 : data_out = 24'b000001101110000011011000;
    16'b0001000000001001 : data_out = 24'b000001101110001010010000;
    16'b0001000000001010 : data_out = 24'b000001101110010001001001;
    16'b0001000000001011 : data_out = 24'b000001101110011000000010;
    16'b0001000000001100 : data_out = 24'b000001101110011110111100;
    16'b0001000000001101 : data_out = 24'b000001101110100101110110;
    16'b0001000000001110 : data_out = 24'b000001101110101100110001;
    16'b0001000000001111 : data_out = 24'b000001101110110011101100;
    16'b0001000000010000 : data_out = 24'b000001101110111010100111;
    16'b0001000000010001 : data_out = 24'b000001101111000001100011;
    16'b0001000000010010 : data_out = 24'b000001101111001000011111;
    16'b0001000000010011 : data_out = 24'b000001101111001111011100;
    16'b0001000000010100 : data_out = 24'b000001101111010110011001;
    16'b0001000000010101 : data_out = 24'b000001101111011101010111;
    16'b0001000000010110 : data_out = 24'b000001101111100100010101;
    16'b0001000000010111 : data_out = 24'b000001101111101011010011;
    16'b0001000000011000 : data_out = 24'b000001101111110010010010;
    16'b0001000000011001 : data_out = 24'b000001101111111001010010;
    16'b0001000000011010 : data_out = 24'b000001110000000000010001;
    16'b0001000000011011 : data_out = 24'b000001110000000111010010;
    16'b0001000000011100 : data_out = 24'b000001110000001110010010;
    16'b0001000000011101 : data_out = 24'b000001110000010101010011;
    16'b0001000000011110 : data_out = 24'b000001110000011100010101;
    16'b0001000000011111 : data_out = 24'b000001110000100011010111;
    16'b0001000000100000 : data_out = 24'b000001110000101010011001;
    16'b0001000000100001 : data_out = 24'b000001110000110001011100;
    16'b0001000000100010 : data_out = 24'b000001110000111000100000;
    16'b0001000000100011 : data_out = 24'b000001110000111111100011;
    16'b0001000000100100 : data_out = 24'b000001110001000110100111;
    16'b0001000000100101 : data_out = 24'b000001110001001101101100;
    16'b0001000000100110 : data_out = 24'b000001110001010100110001;
    16'b0001000000100111 : data_out = 24'b000001110001011011110111;
    16'b0001000000101000 : data_out = 24'b000001110001100010111101;
    16'b0001000000101001 : data_out = 24'b000001110001101010000011;
    16'b0001000000101010 : data_out = 24'b000001110001110001001010;
    16'b0001000000101011 : data_out = 24'b000001110001111000010001;
    16'b0001000000101100 : data_out = 24'b000001110001111111011001;
    16'b0001000000101101 : data_out = 24'b000001110010000110100001;
    16'b0001000000101110 : data_out = 24'b000001110010001101101010;
    16'b0001000000101111 : data_out = 24'b000001110010010100110011;
    16'b0001000000110000 : data_out = 24'b000001110010011011111100;
    16'b0001000000110001 : data_out = 24'b000001110010100011000110;
    16'b0001000000110010 : data_out = 24'b000001110010101010010001;
    16'b0001000000110011 : data_out = 24'b000001110010110001011100;
    16'b0001000000110100 : data_out = 24'b000001110010111000100111;
    16'b0001000000110101 : data_out = 24'b000001110010111111110011;
    16'b0001000000110110 : data_out = 24'b000001110011000110111111;
    16'b0001000000110111 : data_out = 24'b000001110011001110001100;
    16'b0001000000111000 : data_out = 24'b000001110011010101011001;
    16'b0001000000111001 : data_out = 24'b000001110011011100100110;
    16'b0001000000111010 : data_out = 24'b000001110011100011110100;
    16'b0001000000111011 : data_out = 24'b000001110011101011000011;
    16'b0001000000111100 : data_out = 24'b000001110011110010010010;
    16'b0001000000111101 : data_out = 24'b000001110011111001100001;
    16'b0001000000111110 : data_out = 24'b000001110100000000110001;
    16'b0001000000111111 : data_out = 24'b000001110100001000000001;
    16'b0001000001000000 : data_out = 24'b000001110100001111010010;
    16'b0001000001000001 : data_out = 24'b000001110100010110100011;
    16'b0001000001000010 : data_out = 24'b000001110100011101110101;
    16'b0001000001000011 : data_out = 24'b000001110100100101000111;
    16'b0001000001000100 : data_out = 24'b000001110100101100011001;
    16'b0001000001000101 : data_out = 24'b000001110100110011101100;
    16'b0001000001000110 : data_out = 24'b000001110100111011000000;
    16'b0001000001000111 : data_out = 24'b000001110101000010010100;
    16'b0001000001001000 : data_out = 24'b000001110101001001101000;
    16'b0001000001001001 : data_out = 24'b000001110101010000111101;
    16'b0001000001001010 : data_out = 24'b000001110101011000010010;
    16'b0001000001001011 : data_out = 24'b000001110101011111101000;
    16'b0001000001001100 : data_out = 24'b000001110101100110111110;
    16'b0001000001001101 : data_out = 24'b000001110101101110010101;
    16'b0001000001001110 : data_out = 24'b000001110101110101101100;
    16'b0001000001001111 : data_out = 24'b000001110101111101000100;
    16'b0001000001010000 : data_out = 24'b000001110110000100011100;
    16'b0001000001010001 : data_out = 24'b000001110110001011110100;
    16'b0001000001010010 : data_out = 24'b000001110110010011001101;
    16'b0001000001010011 : data_out = 24'b000001110110011010100110;
    16'b0001000001010100 : data_out = 24'b000001110110100010000000;
    16'b0001000001010101 : data_out = 24'b000001110110101001011011;
    16'b0001000001010110 : data_out = 24'b000001110110110000110110;
    16'b0001000001010111 : data_out = 24'b000001110110111000010001;
    16'b0001000001011000 : data_out = 24'b000001110110111111101101;
    16'b0001000001011001 : data_out = 24'b000001110111000111001001;
    16'b0001000001011010 : data_out = 24'b000001110111001110100101;
    16'b0001000001011011 : data_out = 24'b000001110111010110000011;
    16'b0001000001011100 : data_out = 24'b000001110111011101100000;
    16'b0001000001011101 : data_out = 24'b000001110111100100111110;
    16'b0001000001011110 : data_out = 24'b000001110111101100011101;
    16'b0001000001011111 : data_out = 24'b000001110111110011111100;
    16'b0001000001100000 : data_out = 24'b000001110111111011011011;
    16'b0001000001100001 : data_out = 24'b000001111000000010111011;
    16'b0001000001100010 : data_out = 24'b000001111000001010011100;
    16'b0001000001100011 : data_out = 24'b000001111000010001111101;
    16'b0001000001100100 : data_out = 24'b000001111000011001011110;
    16'b0001000001100101 : data_out = 24'b000001111000100001000000;
    16'b0001000001100110 : data_out = 24'b000001111000101000100010;
    16'b0001000001100111 : data_out = 24'b000001111000110000000101;
    16'b0001000001101000 : data_out = 24'b000001111000110111101000;
    16'b0001000001101001 : data_out = 24'b000001111000111111001100;
    16'b0001000001101010 : data_out = 24'b000001111001000110110000;
    16'b0001000001101011 : data_out = 24'b000001111001001110010101;
    16'b0001000001101100 : data_out = 24'b000001111001010101111010;
    16'b0001000001101101 : data_out = 24'b000001111001011101011111;
    16'b0001000001101110 : data_out = 24'b000001111001100101000101;
    16'b0001000001101111 : data_out = 24'b000001111001101100101100;
    16'b0001000001110000 : data_out = 24'b000001111001110100010011;
    16'b0001000001110001 : data_out = 24'b000001111001111011111011;
    16'b0001000001110010 : data_out = 24'b000001111010000011100011;
    16'b0001000001110011 : data_out = 24'b000001111010001011001011;
    16'b0001000001110100 : data_out = 24'b000001111010010010110100;
    16'b0001000001110101 : data_out = 24'b000001111010011010011101;
    16'b0001000001110110 : data_out = 24'b000001111010100010000111;
    16'b0001000001110111 : data_out = 24'b000001111010101001110010;
    16'b0001000001111000 : data_out = 24'b000001111010110001011100;
    16'b0001000001111001 : data_out = 24'b000001111010111001001000;
    16'b0001000001111010 : data_out = 24'b000001111011000000110100;
    16'b0001000001111011 : data_out = 24'b000001111011001000100000;
    16'b0001000001111100 : data_out = 24'b000001111011010000001101;
    16'b0001000001111101 : data_out = 24'b000001111011010111111010;
    16'b0001000001111110 : data_out = 24'b000001111011011111101000;
    16'b0001000001111111 : data_out = 24'b000001111011100111010110;
    16'b0001000010000000 : data_out = 24'b000001111011101111000101;
    16'b0001000010000001 : data_out = 24'b000001111011110110110100;
    16'b0001000010000010 : data_out = 24'b000001111011111110100011;
    16'b0001000010000011 : data_out = 24'b000001111100000110010100;
    16'b0001000010000100 : data_out = 24'b000001111100001110000100;
    16'b0001000010000101 : data_out = 24'b000001111100010101110101;
    16'b0001000010000110 : data_out = 24'b000001111100011101100111;
    16'b0001000010000111 : data_out = 24'b000001111100100101011001;
    16'b0001000010001000 : data_out = 24'b000001111100101101001100;
    16'b0001000010001001 : data_out = 24'b000001111100110100111111;
    16'b0001000010001010 : data_out = 24'b000001111100111100110010;
    16'b0001000010001011 : data_out = 24'b000001111101000100100110;
    16'b0001000010001100 : data_out = 24'b000001111101001100011011;
    16'b0001000010001101 : data_out = 24'b000001111101010100010000;
    16'b0001000010001110 : data_out = 24'b000001111101011100000101;
    16'b0001000010001111 : data_out = 24'b000001111101100011111011;
    16'b0001000010010000 : data_out = 24'b000001111101101011110010;
    16'b0001000010010001 : data_out = 24'b000001111101110011101001;
    16'b0001000010010010 : data_out = 24'b000001111101111011100000;
    16'b0001000010010011 : data_out = 24'b000001111110000011011000;
    16'b0001000010010100 : data_out = 24'b000001111110001011010001;
    16'b0001000010010101 : data_out = 24'b000001111110010011001010;
    16'b0001000010010110 : data_out = 24'b000001111110011011000011;
    16'b0001000010010111 : data_out = 24'b000001111110100010111101;
    16'b0001000010011000 : data_out = 24'b000001111110101010111000;
    16'b0001000010011001 : data_out = 24'b000001111110110010110010;
    16'b0001000010011010 : data_out = 24'b000001111110111010101110;
    16'b0001000010011011 : data_out = 24'b000001111111000010101010;
    16'b0001000010011100 : data_out = 24'b000001111111001010100110;
    16'b0001000010011101 : data_out = 24'b000001111111010010100011;
    16'b0001000010011110 : data_out = 24'b000001111111011010100001;
    16'b0001000010011111 : data_out = 24'b000001111111100010011110;
    16'b0001000010100000 : data_out = 24'b000001111111101010011101;
    16'b0001000010100001 : data_out = 24'b000001111111110010011100;
    16'b0001000010100010 : data_out = 24'b000001111111111010011011;
    16'b0001000010100011 : data_out = 24'b000010000000000010011011;
    16'b0001000010100100 : data_out = 24'b000010000000001010011011;
    16'b0001000010100101 : data_out = 24'b000010000000010010011100;
    16'b0001000010100110 : data_out = 24'b000010000000011010011110;
    16'b0001000010100111 : data_out = 24'b000010000000100010100000;
    16'b0001000010101000 : data_out = 24'b000010000000101010100010;
    16'b0001000010101001 : data_out = 24'b000010000000110010100101;
    16'b0001000010101010 : data_out = 24'b000010000000111010101000;
    16'b0001000010101011 : data_out = 24'b000010000001000010101100;
    16'b0001000010101100 : data_out = 24'b000010000001001010110001;
    16'b0001000010101101 : data_out = 24'b000010000001010010110110;
    16'b0001000010101110 : data_out = 24'b000010000001011010111011;
    16'b0001000010101111 : data_out = 24'b000010000001100011000001;
    16'b0001000010110000 : data_out = 24'b000010000001101011000111;
    16'b0001000010110001 : data_out = 24'b000010000001110011001110;
    16'b0001000010110010 : data_out = 24'b000010000001111011010110;
    16'b0001000010110011 : data_out = 24'b000010000010000011011110;
    16'b0001000010110100 : data_out = 24'b000010000010001011100110;
    16'b0001000010110101 : data_out = 24'b000010000010010011101111;
    16'b0001000010110110 : data_out = 24'b000010000010011011111001;
    16'b0001000010110111 : data_out = 24'b000010000010100100000011;
    16'b0001000010111000 : data_out = 24'b000010000010101100001101;
    16'b0001000010111001 : data_out = 24'b000010000010110100011000;
    16'b0001000010111010 : data_out = 24'b000010000010111100100100;
    16'b0001000010111011 : data_out = 24'b000010000011000100110000;
    16'b0001000010111100 : data_out = 24'b000010000011001100111100;
    16'b0001000010111101 : data_out = 24'b000010000011010101001001;
    16'b0001000010111110 : data_out = 24'b000010000011011101010111;
    16'b0001000010111111 : data_out = 24'b000010000011100101100101;
    16'b0001000011000000 : data_out = 24'b000010000011101101110100;
    16'b0001000011000001 : data_out = 24'b000010000011110110000011;
    16'b0001000011000010 : data_out = 24'b000010000011111110010011;
    16'b0001000011000011 : data_out = 24'b000010000100000110100011;
    16'b0001000011000100 : data_out = 24'b000010000100001110110011;
    16'b0001000011000101 : data_out = 24'b000010000100010111000101;
    16'b0001000011000110 : data_out = 24'b000010000100011111010110;
    16'b0001000011000111 : data_out = 24'b000010000100100111101000;
    16'b0001000011001000 : data_out = 24'b000010000100101111111011;
    16'b0001000011001001 : data_out = 24'b000010000100111000001110;
    16'b0001000011001010 : data_out = 24'b000010000101000000100010;
    16'b0001000011001011 : data_out = 24'b000010000101001000110110;
    16'b0001000011001100 : data_out = 24'b000010000101010001001011;
    16'b0001000011001101 : data_out = 24'b000010000101011001100001;
    16'b0001000011001110 : data_out = 24'b000010000101100001110110;
    16'b0001000011001111 : data_out = 24'b000010000101101010001101;
    16'b0001000011010000 : data_out = 24'b000010000101110010100100;
    16'b0001000011010001 : data_out = 24'b000010000101111010111011;
    16'b0001000011010010 : data_out = 24'b000010000110000011010011;
    16'b0001000011010011 : data_out = 24'b000010000110001011101100;
    16'b0001000011010100 : data_out = 24'b000010000110010100000101;
    16'b0001000011010101 : data_out = 24'b000010000110011100011110;
    16'b0001000011010110 : data_out = 24'b000010000110100100111000;
    16'b0001000011010111 : data_out = 24'b000010000110101101010011;
    16'b0001000011011000 : data_out = 24'b000010000110110101101110;
    16'b0001000011011001 : data_out = 24'b000010000110111110001001;
    16'b0001000011011010 : data_out = 24'b000010000111000110100110;
    16'b0001000011011011 : data_out = 24'b000010000111001111000010;
    16'b0001000011011100 : data_out = 24'b000010000111010111011111;
    16'b0001000011011101 : data_out = 24'b000010000111011111111101;
    16'b0001000011011110 : data_out = 24'b000010000111101000011011;
    16'b0001000011011111 : data_out = 24'b000010000111110000111010;
    16'b0001000011100000 : data_out = 24'b000010000111111001011010;
    16'b0001000011100001 : data_out = 24'b000010001000000001111001;
    16'b0001000011100010 : data_out = 24'b000010001000001010011010;
    16'b0001000011100011 : data_out = 24'b000010001000010010111011;
    16'b0001000011100100 : data_out = 24'b000010001000011011011100;
    16'b0001000011100101 : data_out = 24'b000010001000100011111110;
    16'b0001000011100110 : data_out = 24'b000010001000101100100001;
    16'b0001000011100111 : data_out = 24'b000010001000110101000100;
    16'b0001000011101000 : data_out = 24'b000010001000111101100111;
    16'b0001000011101001 : data_out = 24'b000010001001000110001011;
    16'b0001000011101010 : data_out = 24'b000010001001001110110000;
    16'b0001000011101011 : data_out = 24'b000010001001010111010101;
    16'b0001000011101100 : data_out = 24'b000010001001011111111011;
    16'b0001000011101101 : data_out = 24'b000010001001101000100001;
    16'b0001000011101110 : data_out = 24'b000010001001110001001000;
    16'b0001000011101111 : data_out = 24'b000010001001111001101111;
    16'b0001000011110000 : data_out = 24'b000010001010000010010111;
    16'b0001000011110001 : data_out = 24'b000010001010001011000000;
    16'b0001000011110010 : data_out = 24'b000010001010010011101001;
    16'b0001000011110011 : data_out = 24'b000010001010011100010010;
    16'b0001000011110100 : data_out = 24'b000010001010100100111100;
    16'b0001000011110101 : data_out = 24'b000010001010101101100111;
    16'b0001000011110110 : data_out = 24'b000010001010110110010010;
    16'b0001000011110111 : data_out = 24'b000010001010111110111110;
    16'b0001000011111000 : data_out = 24'b000010001011000111101010;
    16'b0001000011111001 : data_out = 24'b000010001011010000010111;
    16'b0001000011111010 : data_out = 24'b000010001011011001000100;
    16'b0001000011111011 : data_out = 24'b000010001011100001110010;
    16'b0001000011111100 : data_out = 24'b000010001011101010100000;
    16'b0001000011111101 : data_out = 24'b000010001011110011001111;
    16'b0001000011111110 : data_out = 24'b000010001011111011111110;
    16'b0001000011111111 : data_out = 24'b000010001100000100101110;
    16'b0001000100000000 : data_out = 24'b000010001100001101011111;
    16'b0001000100000001 : data_out = 24'b000010001100010110010000;
    16'b0001000100000010 : data_out = 24'b000010001100011111000010;
    16'b0001000100000011 : data_out = 24'b000010001100100111110100;
    16'b0001000100000100 : data_out = 24'b000010001100110000100111;
    16'b0001000100000101 : data_out = 24'b000010001100111001011010;
    16'b0001000100000110 : data_out = 24'b000010001101000010001110;
    16'b0001000100000111 : data_out = 24'b000010001101001011000010;
    16'b0001000100001000 : data_out = 24'b000010001101010011110111;
    16'b0001000100001001 : data_out = 24'b000010001101011100101101;
    16'b0001000100001010 : data_out = 24'b000010001101100101100011;
    16'b0001000100001011 : data_out = 24'b000010001101101110011010;
    16'b0001000100001100 : data_out = 24'b000010001101110111010001;
    16'b0001000100001101 : data_out = 24'b000010001110000000001000;
    16'b0001000100001110 : data_out = 24'b000010001110001001000001;
    16'b0001000100001111 : data_out = 24'b000010001110010001111010;
    16'b0001000100010000 : data_out = 24'b000010001110011010110011;
    16'b0001000100010001 : data_out = 24'b000010001110100011101101;
    16'b0001000100010010 : data_out = 24'b000010001110101100100111;
    16'b0001000100010011 : data_out = 24'b000010001110110101100011;
    16'b0001000100010100 : data_out = 24'b000010001110111110011110;
    16'b0001000100010101 : data_out = 24'b000010001111000111011010;
    16'b0001000100010110 : data_out = 24'b000010001111010000010111;
    16'b0001000100010111 : data_out = 24'b000010001111011001010100;
    16'b0001000100011000 : data_out = 24'b000010001111100010010010;
    16'b0001000100011001 : data_out = 24'b000010001111101011010001;
    16'b0001000100011010 : data_out = 24'b000010001111110100010000;
    16'b0001000100011011 : data_out = 24'b000010001111111101001111;
    16'b0001000100011100 : data_out = 24'b000010010000000110001111;
    16'b0001000100011101 : data_out = 24'b000010010000001111010000;
    16'b0001000100011110 : data_out = 24'b000010010000011000010001;
    16'b0001000100011111 : data_out = 24'b000010010000100001010011;
    16'b0001000100100000 : data_out = 24'b000010010000101010010101;
    16'b0001000100100001 : data_out = 24'b000010010000110011011000;
    16'b0001000100100010 : data_out = 24'b000010010000111100011100;
    16'b0001000100100011 : data_out = 24'b000010010001000101100000;
    16'b0001000100100100 : data_out = 24'b000010010001001110100101;
    16'b0001000100100101 : data_out = 24'b000010010001010111101010;
    16'b0001000100100110 : data_out = 24'b000010010001100000101111;
    16'b0001000100100111 : data_out = 24'b000010010001101001110110;
    16'b0001000100101000 : data_out = 24'b000010010001110010111101;
    16'b0001000100101001 : data_out = 24'b000010010001111100000100;
    16'b0001000100101010 : data_out = 24'b000010010010000101001100;
    16'b0001000100101011 : data_out = 24'b000010010010001110010101;
    16'b0001000100101100 : data_out = 24'b000010010010010111011110;
    16'b0001000100101101 : data_out = 24'b000010010010100000101000;
    16'b0001000100101110 : data_out = 24'b000010010010101001110010;
    16'b0001000100101111 : data_out = 24'b000010010010110010111101;
    16'b0001000100110000 : data_out = 24'b000010010010111100001000;
    16'b0001000100110001 : data_out = 24'b000010010011000101010100;
    16'b0001000100110010 : data_out = 24'b000010010011001110100001;
    16'b0001000100110011 : data_out = 24'b000010010011010111101110;
    16'b0001000100110100 : data_out = 24'b000010010011100000111100;
    16'b0001000100110101 : data_out = 24'b000010010011101010001010;
    16'b0001000100110110 : data_out = 24'b000010010011110011011001;
    16'b0001000100110111 : data_out = 24'b000010010011111100101001;
    16'b0001000100111000 : data_out = 24'b000010010100000101111001;
    16'b0001000100111001 : data_out = 24'b000010010100001111001010;
    16'b0001000100111010 : data_out = 24'b000010010100011000011011;
    16'b0001000100111011 : data_out = 24'b000010010100100001101101;
    16'b0001000100111100 : data_out = 24'b000010010100101010111111;
    16'b0001000100111101 : data_out = 24'b000010010100110100010010;
    16'b0001000100111110 : data_out = 24'b000010010100111101100110;
    16'b0001000100111111 : data_out = 24'b000010010101000110111010;
    16'b0001000101000000 : data_out = 24'b000010010101010000001110;
    16'b0001000101000001 : data_out = 24'b000010010101011001100100;
    16'b0001000101000010 : data_out = 24'b000010010101100010111010;
    16'b0001000101000011 : data_out = 24'b000010010101101100010000;
    16'b0001000101000100 : data_out = 24'b000010010101110101100111;
    16'b0001000101000101 : data_out = 24'b000010010101111110111111;
    16'b0001000101000110 : data_out = 24'b000010010110001000010111;
    16'b0001000101000111 : data_out = 24'b000010010110010001110000;
    16'b0001000101001000 : data_out = 24'b000010010110011011001001;
    16'b0001000101001001 : data_out = 24'b000010010110100100100011;
    16'b0001000101001010 : data_out = 24'b000010010110101101111110;
    16'b0001000101001011 : data_out = 24'b000010010110110111011001;
    16'b0001000101001100 : data_out = 24'b000010010111000000110101;
    16'b0001000101001101 : data_out = 24'b000010010111001010010001;
    16'b0001000101001110 : data_out = 24'b000010010111010011101110;
    16'b0001000101001111 : data_out = 24'b000010010111011101001100;
    16'b0001000101010000 : data_out = 24'b000010010111100110101010;
    16'b0001000101010001 : data_out = 24'b000010010111110000001000;
    16'b0001000101010010 : data_out = 24'b000010010111111001101000;
    16'b0001000101010011 : data_out = 24'b000010011000000011001000;
    16'b0001000101010100 : data_out = 24'b000010011000001100101000;
    16'b0001000101010101 : data_out = 24'b000010011000010110001001;
    16'b0001000101010110 : data_out = 24'b000010011000011111101011;
    16'b0001000101010111 : data_out = 24'b000010011000101001001101;
    16'b0001000101011000 : data_out = 24'b000010011000110010110000;
    16'b0001000101011001 : data_out = 24'b000010011000111100010011;
    16'b0001000101011010 : data_out = 24'b000010011001000101111000;
    16'b0001000101011011 : data_out = 24'b000010011001001111011100;
    16'b0001000101011100 : data_out = 24'b000010011001011001000001;
    16'b0001000101011101 : data_out = 24'b000010011001100010100111;
    16'b0001000101011110 : data_out = 24'b000010011001101100001110;
    16'b0001000101011111 : data_out = 24'b000010011001110101110101;
    16'b0001000101100000 : data_out = 24'b000010011001111111011101;
    16'b0001000101100001 : data_out = 24'b000010011010001001000101;
    16'b0001000101100010 : data_out = 24'b000010011010010010101110;
    16'b0001000101100011 : data_out = 24'b000010011010011100010111;
    16'b0001000101100100 : data_out = 24'b000010011010100110000001;
    16'b0001000101100101 : data_out = 24'b000010011010101111101100;
    16'b0001000101100110 : data_out = 24'b000010011010111001010111;
    16'b0001000101100111 : data_out = 24'b000010011011000011000011;
    16'b0001000101101000 : data_out = 24'b000010011011001100110000;
    16'b0001000101101001 : data_out = 24'b000010011011010110011101;
    16'b0001000101101010 : data_out = 24'b000010011011100000001010;
    16'b0001000101101011 : data_out = 24'b000010011011101001111001;
    16'b0001000101101100 : data_out = 24'b000010011011110011101000;
    16'b0001000101101101 : data_out = 24'b000010011011111101010111;
    16'b0001000101101110 : data_out = 24'b000010011100000111000111;
    16'b0001000101101111 : data_out = 24'b000010011100010000111000;
    16'b0001000101110000 : data_out = 24'b000010011100011010101001;
    16'b0001000101110001 : data_out = 24'b000010011100100100011011;
    16'b0001000101110010 : data_out = 24'b000010011100101110001110;
    16'b0001000101110011 : data_out = 24'b000010011100111000000001;
    16'b0001000101110100 : data_out = 24'b000010011101000001110101;
    16'b0001000101110101 : data_out = 24'b000010011101001011101001;
    16'b0001000101110110 : data_out = 24'b000010011101010101011110;
    16'b0001000101110111 : data_out = 24'b000010011101011111010100;
    16'b0001000101111000 : data_out = 24'b000010011101101001001010;
    16'b0001000101111001 : data_out = 24'b000010011101110011000001;
    16'b0001000101111010 : data_out = 24'b000010011101111100111001;
    16'b0001000101111011 : data_out = 24'b000010011110000110110001;
    16'b0001000101111100 : data_out = 24'b000010011110010000101010;
    16'b0001000101111101 : data_out = 24'b000010011110011010100011;
    16'b0001000101111110 : data_out = 24'b000010011110100100011101;
    16'b0001000101111111 : data_out = 24'b000010011110101110010111;
    16'b0001000110000000 : data_out = 24'b000010011110111000010011;
    16'b0001000110000001 : data_out = 24'b000010011111000010001110;
    16'b0001000110000010 : data_out = 24'b000010011111001100001011;
    16'b0001000110000011 : data_out = 24'b000010011111010110001000;
    16'b0001000110000100 : data_out = 24'b000010011111100000000110;
    16'b0001000110000101 : data_out = 24'b000010011111101010000100;
    16'b0001000110000110 : data_out = 24'b000010011111110100000011;
    16'b0001000110000111 : data_out = 24'b000010011111111110000011;
    16'b0001000110001000 : data_out = 24'b000010100000001000000011;
    16'b0001000110001001 : data_out = 24'b000010100000010010000100;
    16'b0001000110001010 : data_out = 24'b000010100000011100000101;
    16'b0001000110001011 : data_out = 24'b000010100000100110000111;
    16'b0001000110001100 : data_out = 24'b000010100000110000001010;
    16'b0001000110001101 : data_out = 24'b000010100000111010001101;
    16'b0001000110001110 : data_out = 24'b000010100001000100010001;
    16'b0001000110001111 : data_out = 24'b000010100001001110010110;
    16'b0001000110010000 : data_out = 24'b000010100001011000011011;
    16'b0001000110010001 : data_out = 24'b000010100001100010100001;
    16'b0001000110010010 : data_out = 24'b000010100001101100100111;
    16'b0001000110010011 : data_out = 24'b000010100001110110101110;
    16'b0001000110010100 : data_out = 24'b000010100010000000110110;
    16'b0001000110010101 : data_out = 24'b000010100010001010111110;
    16'b0001000110010110 : data_out = 24'b000010100010010101000111;
    16'b0001000110010111 : data_out = 24'b000010100010011111010001;
    16'b0001000110011000 : data_out = 24'b000010100010101001011011;
    16'b0001000110011001 : data_out = 24'b000010100010110011100110;
    16'b0001000110011010 : data_out = 24'b000010100010111101110010;
    16'b0001000110011011 : data_out = 24'b000010100011000111111110;
    16'b0001000110011100 : data_out = 24'b000010100011010010001011;
    16'b0001000110011101 : data_out = 24'b000010100011011100011000;
    16'b0001000110011110 : data_out = 24'b000010100011100110100110;
    16'b0001000110011111 : data_out = 24'b000010100011110000110101;
    16'b0001000110100000 : data_out = 24'b000010100011111011000100;
    16'b0001000110100001 : data_out = 24'b000010100100000101010100;
    16'b0001000110100010 : data_out = 24'b000010100100001111100101;
    16'b0001000110100011 : data_out = 24'b000010100100011001110110;
    16'b0001000110100100 : data_out = 24'b000010100100100100001000;
    16'b0001000110100101 : data_out = 24'b000010100100101110011011;
    16'b0001000110100110 : data_out = 24'b000010100100111000101110;
    16'b0001000110100111 : data_out = 24'b000010100101000011000010;
    16'b0001000110101000 : data_out = 24'b000010100101001101010110;
    16'b0001000110101001 : data_out = 24'b000010100101010111101100;
    16'b0001000110101010 : data_out = 24'b000010100101100010000001;
    16'b0001000110101011 : data_out = 24'b000010100101101100011000;
    16'b0001000110101100 : data_out = 24'b000010100101110110101111;
    16'b0001000110101101 : data_out = 24'b000010100110000001000111;
    16'b0001000110101110 : data_out = 24'b000010100110001011011111;
    16'b0001000110101111 : data_out = 24'b000010100110010101111000;
    16'b0001000110110000 : data_out = 24'b000010100110100000010010;
    16'b0001000110110001 : data_out = 24'b000010100110101010101100;
    16'b0001000110110010 : data_out = 24'b000010100110110101000111;
    16'b0001000110110011 : data_out = 24'b000010100110111111100011;
    16'b0001000110110100 : data_out = 24'b000010100111001001111111;
    16'b0001000110110101 : data_out = 24'b000010100111010100011100;
    16'b0001000110110110 : data_out = 24'b000010100111011110111010;
    16'b0001000110110111 : data_out = 24'b000010100111101001011000;
    16'b0001000110111000 : data_out = 24'b000010100111110011110111;
    16'b0001000110111001 : data_out = 24'b000010100111111110010110;
    16'b0001000110111010 : data_out = 24'b000010101000001000110111;
    16'b0001000110111011 : data_out = 24'b000010101000010011011000;
    16'b0001000110111100 : data_out = 24'b000010101000011101111001;
    16'b0001000110111101 : data_out = 24'b000010101000101000011011;
    16'b0001000110111110 : data_out = 24'b000010101000110010111110;
    16'b0001000110111111 : data_out = 24'b000010101000111101100010;
    16'b0001000111000000 : data_out = 24'b000010101001001000000110;
    16'b0001000111000001 : data_out = 24'b000010101001010010101011;
    16'b0001000111000010 : data_out = 24'b000010101001011101010000;
    16'b0001000111000011 : data_out = 24'b000010101001100111110110;
    16'b0001000111000100 : data_out = 24'b000010101001110010011101;
    16'b0001000111000101 : data_out = 24'b000010101001111101000101;
    16'b0001000111000110 : data_out = 24'b000010101010000111101101;
    16'b0001000111000111 : data_out = 24'b000010101010010010010110;
    16'b0001000111001000 : data_out = 24'b000010101010011100111111;
    16'b0001000111001001 : data_out = 24'b000010101010100111101001;
    16'b0001000111001010 : data_out = 24'b000010101010110010010100;
    16'b0001000111001011 : data_out = 24'b000010101010111100111111;
    16'b0001000111001100 : data_out = 24'b000010101011000111101100;
    16'b0001000111001101 : data_out = 24'b000010101011010010011000;
    16'b0001000111001110 : data_out = 24'b000010101011011101000110;
    16'b0001000111001111 : data_out = 24'b000010101011100111110100;
    16'b0001000111010000 : data_out = 24'b000010101011110010100011;
    16'b0001000111010001 : data_out = 24'b000010101011111101010010;
    16'b0001000111010010 : data_out = 24'b000010101100001000000011;
    16'b0001000111010011 : data_out = 24'b000010101100010010110011;
    16'b0001000111010100 : data_out = 24'b000010101100011101100101;
    16'b0001000111010101 : data_out = 24'b000010101100101000010111;
    16'b0001000111010110 : data_out = 24'b000010101100110011001010;
    16'b0001000111010111 : data_out = 24'b000010101100111101111101;
    16'b0001000111011000 : data_out = 24'b000010101101001000110010;
    16'b0001000111011001 : data_out = 24'b000010101101010011100111;
    16'b0001000111011010 : data_out = 24'b000010101101011110011100;
    16'b0001000111011011 : data_out = 24'b000010101101101001010010;
    16'b0001000111011100 : data_out = 24'b000010101101110100001001;
    16'b0001000111011101 : data_out = 24'b000010101101111111000001;
    16'b0001000111011110 : data_out = 24'b000010101110001001111001;
    16'b0001000111011111 : data_out = 24'b000010101110010100110010;
    16'b0001000111100000 : data_out = 24'b000010101110011111101100;
    16'b0001000111100001 : data_out = 24'b000010101110101010100110;
    16'b0001000111100010 : data_out = 24'b000010101110110101100001;
    16'b0001000111100011 : data_out = 24'b000010101111000000011101;
    16'b0001000111100100 : data_out = 24'b000010101111001011011001;
    16'b0001000111100101 : data_out = 24'b000010101111010110010110;
    16'b0001000111100110 : data_out = 24'b000010101111100001010100;
    16'b0001000111100111 : data_out = 24'b000010101111101100010010;
    16'b0001000111101000 : data_out = 24'b000010101111110111010010;
    16'b0001000111101001 : data_out = 24'b000010110000000010010001;
    16'b0001000111101010 : data_out = 24'b000010110000001101010010;
    16'b0001000111101011 : data_out = 24'b000010110000011000010011;
    16'b0001000111101100 : data_out = 24'b000010110000100011010101;
    16'b0001000111101101 : data_out = 24'b000010110000101110010111;
    16'b0001000111101110 : data_out = 24'b000010110000111001011011;
    16'b0001000111101111 : data_out = 24'b000010110001000100011111;
    16'b0001000111110000 : data_out = 24'b000010110001001111100011;
    16'b0001000111110001 : data_out = 24'b000010110001011010101001;
    16'b0001000111110010 : data_out = 24'b000010110001100101101111;
    16'b0001000111110011 : data_out = 24'b000010110001110000110101;
    16'b0001000111110100 : data_out = 24'b000010110001111011111101;
    16'b0001000111110101 : data_out = 24'b000010110010000111000101;
    16'b0001000111110110 : data_out = 24'b000010110010010010001110;
    16'b0001000111110111 : data_out = 24'b000010110010011101010111;
    16'b0001000111111000 : data_out = 24'b000010110010101000100001;
    16'b0001000111111001 : data_out = 24'b000010110010110011101100;
    16'b0001000111111010 : data_out = 24'b000010110010111110111000;
    16'b0001000111111011 : data_out = 24'b000010110011001010000100;
    16'b0001000111111100 : data_out = 24'b000010110011010101010001;
    16'b0001000111111101 : data_out = 24'b000010110011100000011111;
    16'b0001000111111110 : data_out = 24'b000010110011101011101101;
    16'b0001000111111111 : data_out = 24'b000010110011110110111100;
    16'b0001001000000000 : data_out = 24'b000010110100000010001100;
    16'b0001001000000001 : data_out = 24'b000010110100001101011100;
    16'b0001001000000010 : data_out = 24'b000010110100011000101110;
    16'b0001001000000011 : data_out = 24'b000010110100100011111111;
    16'b0001001000000100 : data_out = 24'b000010110100101111010010;
    16'b0001001000000101 : data_out = 24'b000010110100111010100101;
    16'b0001001000000110 : data_out = 24'b000010110101000101111001;
    16'b0001001000000111 : data_out = 24'b000010110101010001001110;
    16'b0001001000001000 : data_out = 24'b000010110101011100100011;
    16'b0001001000001001 : data_out = 24'b000010110101100111111010;
    16'b0001001000001010 : data_out = 24'b000010110101110011010000;
    16'b0001001000001011 : data_out = 24'b000010110101111110101000;
    16'b0001001000001100 : data_out = 24'b000010110110001010000000;
    16'b0001001000001101 : data_out = 24'b000010110110010101011001;
    16'b0001001000001110 : data_out = 24'b000010110110100000110011;
    16'b0001001000001111 : data_out = 24'b000010110110101100001101;
    16'b0001001000010000 : data_out = 24'b000010110110110111101001;
    16'b0001001000010001 : data_out = 24'b000010110111000011000100;
    16'b0001001000010010 : data_out = 24'b000010110111001110100001;
    16'b0001001000010011 : data_out = 24'b000010110111011001111110;
    16'b0001001000010100 : data_out = 24'b000010110111100101011100;
    16'b0001001000010101 : data_out = 24'b000010110111110000111011;
    16'b0001001000010110 : data_out = 24'b000010110111111100011010;
    16'b0001001000010111 : data_out = 24'b000010111000000111111010;
    16'b0001001000011000 : data_out = 24'b000010111000010011011011;
    16'b0001001000011001 : data_out = 24'b000010111000011110111101;
    16'b0001001000011010 : data_out = 24'b000010111000101010011111;
    16'b0001001000011011 : data_out = 24'b000010111000110110000010;
    16'b0001001000011100 : data_out = 24'b000010111001000001100110;
    16'b0001001000011101 : data_out = 24'b000010111001001101001010;
    16'b0001001000011110 : data_out = 24'b000010111001011000110000;
    16'b0001001000011111 : data_out = 24'b000010111001100100010101;
    16'b0001001000100000 : data_out = 24'b000010111001101111111100;
    16'b0001001000100001 : data_out = 24'b000010111001111011100011;
    16'b0001001000100010 : data_out = 24'b000010111010000111001100;
    16'b0001001000100011 : data_out = 24'b000010111010010010110100;
    16'b0001001000100100 : data_out = 24'b000010111010011110011110;
    16'b0001001000100101 : data_out = 24'b000010111010101010001000;
    16'b0001001000100110 : data_out = 24'b000010111010110101110011;
    16'b0001001000100111 : data_out = 24'b000010111011000001011111;
    16'b0001001000101000 : data_out = 24'b000010111011001101001011;
    16'b0001001000101001 : data_out = 24'b000010111011011000111001;
    16'b0001001000101010 : data_out = 24'b000010111011100100100110;
    16'b0001001000101011 : data_out = 24'b000010111011110000010101;
    16'b0001001000101100 : data_out = 24'b000010111011111100000100;
    16'b0001001000101101 : data_out = 24'b000010111100000111110101;
    16'b0001001000101110 : data_out = 24'b000010111100010011100101;
    16'b0001001000101111 : data_out = 24'b000010111100011111010111;
    16'b0001001000110000 : data_out = 24'b000010111100101011001001;
    16'b0001001000110001 : data_out = 24'b000010111100110110111100;
    16'b0001001000110010 : data_out = 24'b000010111101000010110000;
    16'b0001001000110011 : data_out = 24'b000010111101001110100101;
    16'b0001001000110100 : data_out = 24'b000010111101011010011010;
    16'b0001001000110101 : data_out = 24'b000010111101100110010000;
    16'b0001001000110110 : data_out = 24'b000010111101110010000111;
    16'b0001001000110111 : data_out = 24'b000010111101111101111110;
    16'b0001001000111000 : data_out = 24'b000010111110001001110111;
    16'b0001001000111001 : data_out = 24'b000010111110010101110000;
    16'b0001001000111010 : data_out = 24'b000010111110100001101001;
    16'b0001001000111011 : data_out = 24'b000010111110101101100100;
    16'b0001001000111100 : data_out = 24'b000010111110111001011111;
    16'b0001001000111101 : data_out = 24'b000010111111000101011011;
    16'b0001001000111110 : data_out = 24'b000010111111010001011000;
    16'b0001001000111111 : data_out = 24'b000010111111011101010101;
    16'b0001001001000000 : data_out = 24'b000010111111101001010011;
    16'b0001001001000001 : data_out = 24'b000010111111110101010010;
    16'b0001001001000010 : data_out = 24'b000011000000000001010010;
    16'b0001001001000011 : data_out = 24'b000011000000001101010010;
    16'b0001001001000100 : data_out = 24'b000011000000011001010100;
    16'b0001001001000101 : data_out = 24'b000011000000100101010110;
    16'b0001001001000110 : data_out = 24'b000011000000110001011000;
    16'b0001001001000111 : data_out = 24'b000011000000111101011100;
    16'b0001001001001000 : data_out = 24'b000011000001001001100000;
    16'b0001001001001001 : data_out = 24'b000011000001010101100101;
    16'b0001001001001010 : data_out = 24'b000011000001100001101011;
    16'b0001001001001011 : data_out = 24'b000011000001101101110001;
    16'b0001001001001100 : data_out = 24'b000011000001111001111000;
    16'b0001001001001101 : data_out = 24'b000011000010000110000000;
    16'b0001001001001110 : data_out = 24'b000011000010010010001001;
    16'b0001001001001111 : data_out = 24'b000011000010011110010011;
    16'b0001001001010000 : data_out = 24'b000011000010101010011101;
    16'b0001001001010001 : data_out = 24'b000011000010110110101000;
    16'b0001001001010010 : data_out = 24'b000011000011000010110100;
    16'b0001001001010011 : data_out = 24'b000011000011001111000000;
    16'b0001001001010100 : data_out = 24'b000011000011011011001110;
    16'b0001001001010101 : data_out = 24'b000011000011100111011100;
    16'b0001001001010110 : data_out = 24'b000011000011110011101011;
    16'b0001001001010111 : data_out = 24'b000011000011111111111010;
    16'b0001001001011000 : data_out = 24'b000011000100001100001011;
    16'b0001001001011001 : data_out = 24'b000011000100011000011100;
    16'b0001001001011010 : data_out = 24'b000011000100100100101110;
    16'b0001001001011011 : data_out = 24'b000011000100110001000000;
    16'b0001001001011100 : data_out = 24'b000011000100111101010100;
    16'b0001001001011101 : data_out = 24'b000011000101001001101000;
    16'b0001001001011110 : data_out = 24'b000011000101010101111101;
    16'b0001001001011111 : data_out = 24'b000011000101100010010011;
    16'b0001001001100000 : data_out = 24'b000011000101101110101001;
    16'b0001001001100001 : data_out = 24'b000011000101111011000001;
    16'b0001001001100010 : data_out = 24'b000011000110000111011001;
    16'b0001001001100011 : data_out = 24'b000011000110010011110010;
    16'b0001001001100100 : data_out = 24'b000011000110100000001011;
    16'b0001001001100101 : data_out = 24'b000011000110101100100110;
    16'b0001001001100110 : data_out = 24'b000011000110111001000001;
    16'b0001001001100111 : data_out = 24'b000011000111000101011101;
    16'b0001001001101000 : data_out = 24'b000011000111010001111001;
    16'b0001001001101001 : data_out = 24'b000011000111011110010111;
    16'b0001001001101010 : data_out = 24'b000011000111101010110101;
    16'b0001001001101011 : data_out = 24'b000011000111110111010100;
    16'b0001001001101100 : data_out = 24'b000011001000000011110100;
    16'b0001001001101101 : data_out = 24'b000011001000010000010101;
    16'b0001001001101110 : data_out = 24'b000011001000011100110110;
    16'b0001001001101111 : data_out = 24'b000011001000101001011000;
    16'b0001001001110000 : data_out = 24'b000011001000110101111011;
    16'b0001001001110001 : data_out = 24'b000011001001000010011111;
    16'b0001001001110010 : data_out = 24'b000011001001001111000100;
    16'b0001001001110011 : data_out = 24'b000011001001011011101001;
    16'b0001001001110100 : data_out = 24'b000011001001101000001111;
    16'b0001001001110101 : data_out = 24'b000011001001110100110110;
    16'b0001001001110110 : data_out = 24'b000011001010000001011110;
    16'b0001001001110111 : data_out = 24'b000011001010001110000110;
    16'b0001001001111000 : data_out = 24'b000011001010011010101111;
    16'b0001001001111001 : data_out = 24'b000011001010100111011010;
    16'b0001001001111010 : data_out = 24'b000011001010110100000100;
    16'b0001001001111011 : data_out = 24'b000011001011000000110000;
    16'b0001001001111100 : data_out = 24'b000011001011001101011100;
    16'b0001001001111101 : data_out = 24'b000011001011011010001010;
    16'b0001001001111110 : data_out = 24'b000011001011100110111000;
    16'b0001001001111111 : data_out = 24'b000011001011110011100111;
    16'b0001001010000000 : data_out = 24'b000011001100000000010110;
    16'b0001001010000001 : data_out = 24'b000011001100001101000111;
    16'b0001001010000010 : data_out = 24'b000011001100011001111000;
    16'b0001001010000011 : data_out = 24'b000011001100100110101010;
    16'b0001001010000100 : data_out = 24'b000011001100110011011101;
    16'b0001001010000101 : data_out = 24'b000011001101000000010000;
    16'b0001001010000110 : data_out = 24'b000011001101001101000101;
    16'b0001001010000111 : data_out = 24'b000011001101011001111010;
    16'b0001001010001000 : data_out = 24'b000011001101100110110000;
    16'b0001001010001001 : data_out = 24'b000011001101110011100111;
    16'b0001001010001010 : data_out = 24'b000011001110000000011110;
    16'b0001001010001011 : data_out = 24'b000011001110001101010111;
    16'b0001001010001100 : data_out = 24'b000011001110011010010000;
    16'b0001001010001101 : data_out = 24'b000011001110100111001010;
    16'b0001001010001110 : data_out = 24'b000011001110110100000101;
    16'b0001001010001111 : data_out = 24'b000011001111000001000001;
    16'b0001001010010000 : data_out = 24'b000011001111001101111101;
    16'b0001001010010001 : data_out = 24'b000011001111011010111010;
    16'b0001001010010010 : data_out = 24'b000011001111100111111000;
    16'b0001001010010011 : data_out = 24'b000011001111110100110111;
    16'b0001001010010100 : data_out = 24'b000011010000000001110111;
    16'b0001001010010101 : data_out = 24'b000011010000001110111000;
    16'b0001001010010110 : data_out = 24'b000011010000011011111001;
    16'b0001001010010111 : data_out = 24'b000011010000101000111011;
    16'b0001001010011000 : data_out = 24'b000011010000110101111110;
    16'b0001001010011001 : data_out = 24'b000011010001000011000010;
    16'b0001001010011010 : data_out = 24'b000011010001010000000110;
    16'b0001001010011011 : data_out = 24'b000011010001011101001100;
    16'b0001001010011100 : data_out = 24'b000011010001101010010010;
    16'b0001001010011101 : data_out = 24'b000011010001110111011001;
    16'b0001001010011110 : data_out = 24'b000011010010000100100001;
    16'b0001001010011111 : data_out = 24'b000011010010010001101010;
    16'b0001001010100000 : data_out = 24'b000011010010011110110011;
    16'b0001001010100001 : data_out = 24'b000011010010101011111110;
    16'b0001001010100010 : data_out = 24'b000011010010111001001001;
    16'b0001001010100011 : data_out = 24'b000011010011000110010101;
    16'b0001001010100100 : data_out = 24'b000011010011010011100010;
    16'b0001001010100101 : data_out = 24'b000011010011100000101111;
    16'b0001001010100110 : data_out = 24'b000011010011101101111110;
    16'b0001001010100111 : data_out = 24'b000011010011111011001101;
    16'b0001001010101000 : data_out = 24'b000011010100001000011101;
    16'b0001001010101001 : data_out = 24'b000011010100010101101110;
    16'b0001001010101010 : data_out = 24'b000011010100100011000000;
    16'b0001001010101011 : data_out = 24'b000011010100110000010010;
    16'b0001001010101100 : data_out = 24'b000011010100111101100110;
    16'b0001001010101101 : data_out = 24'b000011010101001010111010;
    16'b0001001010101110 : data_out = 24'b000011010101011000001111;
    16'b0001001010101111 : data_out = 24'b000011010101100101100101;
    16'b0001001010110000 : data_out = 24'b000011010101110010111100;
    16'b0001001010110001 : data_out = 24'b000011010110000000010011;
    16'b0001001010110010 : data_out = 24'b000011010110001101101100;
    16'b0001001010110011 : data_out = 24'b000011010110011011000101;
    16'b0001001010110100 : data_out = 24'b000011010110101000011111;
    16'b0001001010110101 : data_out = 24'b000011010110110101111010;
    16'b0001001010110110 : data_out = 24'b000011010111000011010110;
    16'b0001001010110111 : data_out = 24'b000011010111010000110011;
    16'b0001001010111000 : data_out = 24'b000011010111011110010000;
    16'b0001001010111001 : data_out = 24'b000011010111101011101110;
    16'b0001001010111010 : data_out = 24'b000011010111111001001110;
    16'b0001001010111011 : data_out = 24'b000011011000000110101110;
    16'b0001001010111100 : data_out = 24'b000011011000010100001110;
    16'b0001001010111101 : data_out = 24'b000011011000100001110000;
    16'b0001001010111110 : data_out = 24'b000011011000101111010011;
    16'b0001001010111111 : data_out = 24'b000011011000111100110110;
    16'b0001001011000000 : data_out = 24'b000011011001001010011010;
    16'b0001001011000001 : data_out = 24'b000011011001010111111111;
    16'b0001001011000010 : data_out = 24'b000011011001100101100101;
    16'b0001001011000011 : data_out = 24'b000011011001110011001100;
    16'b0001001011000100 : data_out = 24'b000011011010000000110100;
    16'b0001001011000101 : data_out = 24'b000011011010001110011100;
    16'b0001001011000110 : data_out = 24'b000011011010011100000101;
    16'b0001001011000111 : data_out = 24'b000011011010101001110000;
    16'b0001001011001000 : data_out = 24'b000011011010110111011011;
    16'b0001001011001001 : data_out = 24'b000011011011000101000111;
    16'b0001001011001010 : data_out = 24'b000011011011010010110011;
    16'b0001001011001011 : data_out = 24'b000011011011100000100001;
    16'b0001001011001100 : data_out = 24'b000011011011101110001111;
    16'b0001001011001101 : data_out = 24'b000011011011111011111111;
    16'b0001001011001110 : data_out = 24'b000011011100001001101111;
    16'b0001001011001111 : data_out = 24'b000011011100010111100000;
    16'b0001001011010000 : data_out = 24'b000011011100100101010010;
    16'b0001001011010001 : data_out = 24'b000011011100110011000101;
    16'b0001001011010010 : data_out = 24'b000011011101000000111000;
    16'b0001001011010011 : data_out = 24'b000011011101001110101101;
    16'b0001001011010100 : data_out = 24'b000011011101011100100010;
    16'b0001001011010101 : data_out = 24'b000011011101101010011000;
    16'b0001001011010110 : data_out = 24'b000011011101111000001111;
    16'b0001001011010111 : data_out = 24'b000011011110000110000111;
    16'b0001001011011000 : data_out = 24'b000011011110010100000000;
    16'b0001001011011001 : data_out = 24'b000011011110100001111010;
    16'b0001001011011010 : data_out = 24'b000011011110101111110100;
    16'b0001001011011011 : data_out = 24'b000011011110111101110000;
    16'b0001001011011100 : data_out = 24'b000011011111001011101100;
    16'b0001001011011101 : data_out = 24'b000011011111011001101001;
    16'b0001001011011110 : data_out = 24'b000011011111100111100111;
    16'b0001001011011111 : data_out = 24'b000011011111110101100110;
    16'b0001001011100000 : data_out = 24'b000011100000000011100110;
    16'b0001001011100001 : data_out = 24'b000011100000010001100111;
    16'b0001001011100010 : data_out = 24'b000011100000011111101000;
    16'b0001001011100011 : data_out = 24'b000011100000101101101011;
    16'b0001001011100100 : data_out = 24'b000011100000111011101110;
    16'b0001001011100101 : data_out = 24'b000011100001001001110010;
    16'b0001001011100110 : data_out = 24'b000011100001010111110111;
    16'b0001001011100111 : data_out = 24'b000011100001100101111101;
    16'b0001001011101000 : data_out = 24'b000011100001110100000100;
    16'b0001001011101001 : data_out = 24'b000011100010000010001100;
    16'b0001001011101010 : data_out = 24'b000011100010010000010100;
    16'b0001001011101011 : data_out = 24'b000011100010011110011110;
    16'b0001001011101100 : data_out = 24'b000011100010101100101000;
    16'b0001001011101101 : data_out = 24'b000011100010111010110011;
    16'b0001001011101110 : data_out = 24'b000011100011001000111111;
    16'b0001001011101111 : data_out = 24'b000011100011010111001100;
    16'b0001001011110000 : data_out = 24'b000011100011100101011010;
    16'b0001001011110001 : data_out = 24'b000011100011110011101001;
    16'b0001001011110010 : data_out = 24'b000011100100000001111001;
    16'b0001001011110011 : data_out = 24'b000011100100010000001001;
    16'b0001001011110100 : data_out = 24'b000011100100011110011011;
    16'b0001001011110101 : data_out = 24'b000011100100101100101101;
    16'b0001001011110110 : data_out = 24'b000011100100111011000000;
    16'b0001001011110111 : data_out = 24'b000011100101001001010100;
    16'b0001001011111000 : data_out = 24'b000011100101010111101001;
    16'b0001001011111001 : data_out = 24'b000011100101100101111111;
    16'b0001001011111010 : data_out = 24'b000011100101110100010110;
    16'b0001001011111011 : data_out = 24'b000011100110000010101110;
    16'b0001001011111100 : data_out = 24'b000011100110010001000110;
    16'b0001001011111101 : data_out = 24'b000011100110011111100000;
    16'b0001001011111110 : data_out = 24'b000011100110101101111010;
    16'b0001001011111111 : data_out = 24'b000011100110111100010110;
    16'b0001001100000000 : data_out = 24'b000011100111001010110010;
    16'b0001001100000001 : data_out = 24'b000011100111011001001111;
    16'b0001001100000010 : data_out = 24'b000011100111100111101101;
    16'b0001001100000011 : data_out = 24'b000011100111110110001100;
    16'b0001001100000100 : data_out = 24'b000011101000000100101100;
    16'b0001001100000101 : data_out = 24'b000011101000010011001101;
    16'b0001001100000110 : data_out = 24'b000011101000100001101110;
    16'b0001001100000111 : data_out = 24'b000011101000110000010001;
    16'b0001001100001000 : data_out = 24'b000011101000111110110100;
    16'b0001001100001001 : data_out = 24'b000011101001001101011001;
    16'b0001001100001010 : data_out = 24'b000011101001011011111110;
    16'b0001001100001011 : data_out = 24'b000011101001101010100100;
    16'b0001001100001100 : data_out = 24'b000011101001111001001011;
    16'b0001001100001101 : data_out = 24'b000011101010000111110011;
    16'b0001001100001110 : data_out = 24'b000011101010010110011100;
    16'b0001001100001111 : data_out = 24'b000011101010100101000110;
    16'b0001001100010000 : data_out = 24'b000011101010110011110001;
    16'b0001001100010001 : data_out = 24'b000011101011000010011101;
    16'b0001001100010010 : data_out = 24'b000011101011010001001001;
    16'b0001001100010011 : data_out = 24'b000011101011011111110111;
    16'b0001001100010100 : data_out = 24'b000011101011101110100101;
    16'b0001001100010101 : data_out = 24'b000011101011111101010101;
    16'b0001001100010110 : data_out = 24'b000011101100001100000101;
    16'b0001001100010111 : data_out = 24'b000011101100011010110110;
    16'b0001001100011000 : data_out = 24'b000011101100101001101000;
    16'b0001001100011001 : data_out = 24'b000011101100111000011011;
    16'b0001001100011010 : data_out = 24'b000011101101000111001111;
    16'b0001001100011011 : data_out = 24'b000011101101010110000100;
    16'b0001001100011100 : data_out = 24'b000011101101100100111010;
    16'b0001001100011101 : data_out = 24'b000011101101110011110001;
    16'b0001001100011110 : data_out = 24'b000011101110000010101001;
    16'b0001001100011111 : data_out = 24'b000011101110010001100001;
    16'b0001001100100000 : data_out = 24'b000011101110100000011011;
    16'b0001001100100001 : data_out = 24'b000011101110101111010101;
    16'b0001001100100010 : data_out = 24'b000011101110111110010001;
    16'b0001001100100011 : data_out = 24'b000011101111001101001101;
    16'b0001001100100100 : data_out = 24'b000011101111011100001010;
    16'b0001001100100101 : data_out = 24'b000011101111101011001001;
    16'b0001001100100110 : data_out = 24'b000011101111111010001000;
    16'b0001001100100111 : data_out = 24'b000011110000001001001000;
    16'b0001001100101000 : data_out = 24'b000011110000011000001001;
    16'b0001001100101001 : data_out = 24'b000011110000100111001011;
    16'b0001001100101010 : data_out = 24'b000011110000110110001110;
    16'b0001001100101011 : data_out = 24'b000011110001000101010010;
    16'b0001001100101100 : data_out = 24'b000011110001010100010110;
    16'b0001001100101101 : data_out = 24'b000011110001100011011100;
    16'b0001001100101110 : data_out = 24'b000011110001110010100011;
    16'b0001001100101111 : data_out = 24'b000011110010000001101010;
    16'b0001001100110000 : data_out = 24'b000011110010010000110011;
    16'b0001001100110001 : data_out = 24'b000011110010011111111101;
    16'b0001001100110010 : data_out = 24'b000011110010101111000111;
    16'b0001001100110011 : data_out = 24'b000011110010111110010010;
    16'b0001001100110100 : data_out = 24'b000011110011001101011111;
    16'b0001001100110101 : data_out = 24'b000011110011011100101100;
    16'b0001001100110110 : data_out = 24'b000011110011101011111010;
    16'b0001001100110111 : data_out = 24'b000011110011111011001010;
    16'b0001001100111000 : data_out = 24'b000011110100001010011010;
    16'b0001001100111001 : data_out = 24'b000011110100011001101011;
    16'b0001001100111010 : data_out = 24'b000011110100101000111101;
    16'b0001001100111011 : data_out = 24'b000011110100111000010000;
    16'b0001001100111100 : data_out = 24'b000011110101000111100100;
    16'b0001001100111101 : data_out = 24'b000011110101010110111001;
    16'b0001001100111110 : data_out = 24'b000011110101100110001111;
    16'b0001001100111111 : data_out = 24'b000011110101110101100110;
    16'b0001001101000000 : data_out = 24'b000011110110000100111110;
    16'b0001001101000001 : data_out = 24'b000011110110010100010110;
    16'b0001001101000010 : data_out = 24'b000011110110100011110000;
    16'b0001001101000011 : data_out = 24'b000011110110110011001011;
    16'b0001001101000100 : data_out = 24'b000011110111000010100111;
    16'b0001001101000101 : data_out = 24'b000011110111010010000011;
    16'b0001001101000110 : data_out = 24'b000011110111100001100001;
    16'b0001001101000111 : data_out = 24'b000011110111110000111111;
    16'b0001001101001000 : data_out = 24'b000011111000000000011111;
    16'b0001001101001001 : data_out = 24'b000011111000001111111111;
    16'b0001001101001010 : data_out = 24'b000011111000011111100001;
    16'b0001001101001011 : data_out = 24'b000011111000101111000011;
    16'b0001001101001100 : data_out = 24'b000011111000111110100111;
    16'b0001001101001101 : data_out = 24'b000011111001001110001011;
    16'b0001001101001110 : data_out = 24'b000011111001011101110001;
    16'b0001001101001111 : data_out = 24'b000011111001101101010111;
    16'b0001001101010000 : data_out = 24'b000011111001111100111110;
    16'b0001001101010001 : data_out = 24'b000011111010001100100111;
    16'b0001001101010010 : data_out = 24'b000011111010011100010000;
    16'b0001001101010011 : data_out = 24'b000011111010101011111010;
    16'b0001001101010100 : data_out = 24'b000011111010111011100101;
    16'b0001001101010101 : data_out = 24'b000011111011001011010010;
    16'b0001001101010110 : data_out = 24'b000011111011011010111111;
    16'b0001001101010111 : data_out = 24'b000011111011101010101101;
    16'b0001001101011000 : data_out = 24'b000011111011111010011100;
    16'b0001001101011001 : data_out = 24'b000011111100001010001100;
    16'b0001001101011010 : data_out = 24'b000011111100011001111101;
    16'b0001001101011011 : data_out = 24'b000011111100101001101111;
    16'b0001001101011100 : data_out = 24'b000011111100111001100011;
    16'b0001001101011101 : data_out = 24'b000011111101001001010111;
    16'b0001001101011110 : data_out = 24'b000011111101011001001100;
    16'b0001001101011111 : data_out = 24'b000011111101101001000010;
    16'b0001001101100000 : data_out = 24'b000011111101111000111001;
    16'b0001001101100001 : data_out = 24'b000011111110001000110001;
    16'b0001001101100010 : data_out = 24'b000011111110011000101010;
    16'b0001001101100011 : data_out = 24'b000011111110101000100100;
    16'b0001001101100100 : data_out = 24'b000011111110111000011111;
    16'b0001001101100101 : data_out = 24'b000011111111001000011011;
    16'b0001001101100110 : data_out = 24'b000011111111011000011000;
    16'b0001001101100111 : data_out = 24'b000011111111101000010110;
    16'b0001001101101000 : data_out = 24'b000011111111111000010101;
    16'b0001001101101001 : data_out = 24'b000100000000001000010101;
    16'b0001001101101010 : data_out = 24'b000100000000011000010110;
    16'b0001001101101011 : data_out = 24'b000100000000101000011000;
    16'b0001001101101100 : data_out = 24'b000100000000111000011011;
    16'b0001001101101101 : data_out = 24'b000100000001001000011111;
    16'b0001001101101110 : data_out = 24'b000100000001011000100100;
    16'b0001001101101111 : data_out = 24'b000100000001101000101010;
    16'b0001001101110000 : data_out = 24'b000100000001111000110001;
    16'b0001001101110001 : data_out = 24'b000100000010001000111001;
    16'b0001001101110010 : data_out = 24'b000100000010011001000010;
    16'b0001001101110011 : data_out = 24'b000100000010101001001101;
    16'b0001001101110100 : data_out = 24'b000100000010111001011000;
    16'b0001001101110101 : data_out = 24'b000100000011001001100100;
    16'b0001001101110110 : data_out = 24'b000100000011011001110001;
    16'b0001001101110111 : data_out = 24'b000100000011101001111111;
    16'b0001001101111000 : data_out = 24'b000100000011111010001110;
    16'b0001001101111001 : data_out = 24'b000100000100001010011110;
    16'b0001001101111010 : data_out = 24'b000100000100011010101111;
    16'b0001001101111011 : data_out = 24'b000100000100101011000010;
    16'b0001001101111100 : data_out = 24'b000100000100111011010101;
    16'b0001001101111101 : data_out = 24'b000100000101001011101001;
    16'b0001001101111110 : data_out = 24'b000100000101011011111110;
    16'b0001001101111111 : data_out = 24'b000100000101101100010100;
    16'b0001001110000000 : data_out = 24'b000100000101111100101100;
    16'b0001001110000001 : data_out = 24'b000100000110001101000100;
    16'b0001001110000010 : data_out = 24'b000100000110011101011101;
    16'b0001001110000011 : data_out = 24'b000100000110101101111000;
    16'b0001001110000100 : data_out = 24'b000100000110111110010011;
    16'b0001001110000101 : data_out = 24'b000100000111001110110000;
    16'b0001001110000110 : data_out = 24'b000100000111011111001101;
    16'b0001001110000111 : data_out = 24'b000100000111101111101011;
    16'b0001001110001000 : data_out = 24'b000100001000000000001011;
    16'b0001001110001001 : data_out = 24'b000100001000010000101011;
    16'b0001001110001010 : data_out = 24'b000100001000100001001101;
    16'b0001001110001011 : data_out = 24'b000100001000110001110000;
    16'b0001001110001100 : data_out = 24'b000100001001000010010011;
    16'b0001001110001101 : data_out = 24'b000100001001010010111000;
    16'b0001001110001110 : data_out = 24'b000100001001100011011110;
    16'b0001001110001111 : data_out = 24'b000100001001110100000100;
    16'b0001001110010000 : data_out = 24'b000100001010000100101100;
    16'b0001001110010001 : data_out = 24'b000100001010010101010101;
    16'b0001001110010010 : data_out = 24'b000100001010100101111111;
    16'b0001001110010011 : data_out = 24'b000100001010110110101010;
    16'b0001001110010100 : data_out = 24'b000100001011000111010110;
    16'b0001001110010101 : data_out = 24'b000100001011011000000011;
    16'b0001001110010110 : data_out = 24'b000100001011101000110001;
    16'b0001001110010111 : data_out = 24'b000100001011111001100000;
    16'b0001001110011000 : data_out = 24'b000100001100001010010000;
    16'b0001001110011001 : data_out = 24'b000100001100011011000001;
    16'b0001001110011010 : data_out = 24'b000100001100101011110011;
    16'b0001001110011011 : data_out = 24'b000100001100111100100110;
    16'b0001001110011100 : data_out = 24'b000100001101001101011011;
    16'b0001001110011101 : data_out = 24'b000100001101011110010000;
    16'b0001001110011110 : data_out = 24'b000100001101101111000111;
    16'b0001001110011111 : data_out = 24'b000100001101111111111110;
    16'b0001001110100000 : data_out = 24'b000100001110010000110111;
    16'b0001001110100001 : data_out = 24'b000100001110100001110000;
    16'b0001001110100010 : data_out = 24'b000100001110110010101011;
    16'b0001001110100011 : data_out = 24'b000100001111000011100110;
    16'b0001001110100100 : data_out = 24'b000100001111010100100011;
    16'b0001001110100101 : data_out = 24'b000100001111100101100001;
    16'b0001001110100110 : data_out = 24'b000100001111110110100000;
    16'b0001001110100111 : data_out = 24'b000100010000000111100000;
    16'b0001001110101000 : data_out = 24'b000100010000011000100001;
    16'b0001001110101001 : data_out = 24'b000100010000101001100011;
    16'b0001001110101010 : data_out = 24'b000100010000111010100110;
    16'b0001001110101011 : data_out = 24'b000100010001001011101010;
    16'b0001001110101100 : data_out = 24'b000100010001011100101111;
    16'b0001001110101101 : data_out = 24'b000100010001101101110110;
    16'b0001001110101110 : data_out = 24'b000100010001111110111101;
    16'b0001001110101111 : data_out = 24'b000100010010010000000110;
    16'b0001001110110000 : data_out = 24'b000100010010100001001111;
    16'b0001001110110001 : data_out = 24'b000100010010110010011010;
    16'b0001001110110010 : data_out = 24'b000100010011000011100110;
    16'b0001001110110011 : data_out = 24'b000100010011010100110010;
    16'b0001001110110100 : data_out = 24'b000100010011100110000000;
    16'b0001001110110101 : data_out = 24'b000100010011110111001111;
    16'b0001001110110110 : data_out = 24'b000100010100001000011111;
    16'b0001001110110111 : data_out = 24'b000100010100011001110000;
    16'b0001001110111000 : data_out = 24'b000100010100101011000010;
    16'b0001001110111001 : data_out = 24'b000100010100111100010101;
    16'b0001001110111010 : data_out = 24'b000100010101001101101010;
    16'b0001001110111011 : data_out = 24'b000100010101011110111111;
    16'b0001001110111100 : data_out = 24'b000100010101110000010110;
    16'b0001001110111101 : data_out = 24'b000100010110000001101101;
    16'b0001001110111110 : data_out = 24'b000100010110010011000110;
    16'b0001001110111111 : data_out = 24'b000100010110100100100000;
    16'b0001001111000000 : data_out = 24'b000100010110110101111010;
    16'b0001001111000001 : data_out = 24'b000100010111000111010110;
    16'b0001001111000010 : data_out = 24'b000100010111011000110011;
    16'b0001001111000011 : data_out = 24'b000100010111101010010001;
    16'b0001001111000100 : data_out = 24'b000100010111111011110001;
    16'b0001001111000101 : data_out = 24'b000100011000001101010001;
    16'b0001001111000110 : data_out = 24'b000100011000011110110010;
    16'b0001001111000111 : data_out = 24'b000100011000110000010101;
    16'b0001001111001000 : data_out = 24'b000100011001000001111000;
    16'b0001001111001001 : data_out = 24'b000100011001010011011101;
    16'b0001001111001010 : data_out = 24'b000100011001100101000011;
    16'b0001001111001011 : data_out = 24'b000100011001110110101010;
    16'b0001001111001100 : data_out = 24'b000100011010001000010010;
    16'b0001001111001101 : data_out = 24'b000100011010011001111011;
    16'b0001001111001110 : data_out = 24'b000100011010101011100101;
    16'b0001001111001111 : data_out = 24'b000100011010111101010000;
    16'b0001001111010000 : data_out = 24'b000100011011001110111101;
    16'b0001001111010001 : data_out = 24'b000100011011100000101010;
    16'b0001001111010010 : data_out = 24'b000100011011110010011001;
    16'b0001001111010011 : data_out = 24'b000100011100000100001000;
    16'b0001001111010100 : data_out = 24'b000100011100010101111001;
    16'b0001001111010101 : data_out = 24'b000100011100100111101011;
    16'b0001001111010110 : data_out = 24'b000100011100111001011110;
    16'b0001001111010111 : data_out = 24'b000100011101001011010010;
    16'b0001001111011000 : data_out = 24'b000100011101011101001000;
    16'b0001001111011001 : data_out = 24'b000100011101101110111110;
    16'b0001001111011010 : data_out = 24'b000100011110000000110101;
    16'b0001001111011011 : data_out = 24'b000100011110010010101110;
    16'b0001001111011100 : data_out = 24'b000100011110100100101000;
    16'b0001001111011101 : data_out = 24'b000100011110110110100011;
    16'b0001001111011110 : data_out = 24'b000100011111001000011111;
    16'b0001001111011111 : data_out = 24'b000100011111011010011100;
    16'b0001001111100000 : data_out = 24'b000100011111101100011010;
    16'b0001001111100001 : data_out = 24'b000100011111111110011001;
    16'b0001001111100010 : data_out = 24'b000100100000010000011010;
    16'b0001001111100011 : data_out = 24'b000100100000100010011011;
    16'b0001001111100100 : data_out = 24'b000100100000110100011110;
    16'b0001001111100101 : data_out = 24'b000100100001000110100010;
    16'b0001001111100110 : data_out = 24'b000100100001011000100111;
    16'b0001001111100111 : data_out = 24'b000100100001101010101101;
    16'b0001001111101000 : data_out = 24'b000100100001111100110100;
    16'b0001001111101001 : data_out = 24'b000100100010001110111100;
    16'b0001001111101010 : data_out = 24'b000100100010100001000110;
    16'b0001001111101011 : data_out = 24'b000100100010110011010001;
    16'b0001001111101100 : data_out = 24'b000100100011000101011100;
    16'b0001001111101101 : data_out = 24'b000100100011010111101001;
    16'b0001001111101110 : data_out = 24'b000100100011101001110111;
    16'b0001001111101111 : data_out = 24'b000100100011111100000111;
    16'b0001001111110000 : data_out = 24'b000100100100001110010111;
    16'b0001001111110001 : data_out = 24'b000100100100100000101000;
    16'b0001001111110010 : data_out = 24'b000100100100110010111011;
    16'b0001001111110011 : data_out = 24'b000100100101000101001111;
    16'b0001001111110100 : data_out = 24'b000100100101010111100100;
    16'b0001001111110101 : data_out = 24'b000100100101101001111010;
    16'b0001001111110110 : data_out = 24'b000100100101111100010001;
    16'b0001001111110111 : data_out = 24'b000100100110001110101001;
    16'b0001001111111000 : data_out = 24'b000100100110100001000011;
    16'b0001001111111001 : data_out = 24'b000100100110110011011101;
    16'b0001001111111010 : data_out = 24'b000100100111000101111001;
    16'b0001001111111011 : data_out = 24'b000100100111011000010110;
    16'b0001001111111100 : data_out = 24'b000100100111101010110100;
    16'b0001001111111101 : data_out = 24'b000100100111111101010011;
    16'b0001001111111110 : data_out = 24'b000100101000001111110100;
    16'b0001001111111111 : data_out = 24'b000100101000100010010101;
    16'b0001010000000000 : data_out = 24'b000100101000110100111000;
	endcase
end
endmodule

