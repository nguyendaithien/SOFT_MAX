module LUT #(parameter DATA_WIDTH = 16 , DATA_WIDTH_OUT = 24) (
		data_in
	 ,data_out
);
	input [DATA_WIDTH-1:0] data_in;
	output reg [DATA_WIDTH_OUT-1:0] data_out;
always @(data_in) begin
	case(data_in) 	
		16'b1101100000000000 : data_out =  24'b000000000000000000011011;
		16'b1101100000000011 : data_out =  24'b000000000000000000011011;
		16'b1101100000000101 : data_out =  24'b000000000000000000011011;
		16'b1101100000000111 : data_out =  24'b000000000000000000011011;
		16'b1101100000001001 : data_out =  24'b000000000000000000011011;
		16'b1101100000001011 : data_out =  24'b000000000000000000011011;
		16'b1101100000001101 : data_out =  24'b000000000000000000011011;
		16'b1101100000001111 : data_out =  24'b000000000000000000011011;
		16'b1101100000010001 : data_out =  24'b000000000000000000011011;
		16'b1101100000010011 : data_out =  24'b000000000000000000011011;
		16'b1101100000010101 : data_out =  24'b000000000000000000011011;
		16'b1101100000010111 : data_out =  24'b000000000000000000011011;
		16'b1101100000011001 : data_out =  24'b000000000000000000011011;
		16'b1101100000011011 : data_out =  24'b000000000000000000011011;
		16'b1101100000011101 : data_out =  24'b000000000000000000011011;
		16'b1101100000011111 : data_out =  24'b000000000000000000011100;
		16'b1101100000100001 : data_out =  24'b000000000000000000011100;
		16'b1101100000100011 : data_out =  24'b000000000000000000011100;
		16'b1101100000100101 : data_out =  24'b000000000000000000011100;
		16'b1101100000100111 : data_out =  24'b000000000000000000011100;
		16'b1101100000101001 : data_out =  24'b000000000000000000011100;
		16'b1101100000101100 : data_out =  24'b000000000000000000011100;
		16'b1101100000101110 : data_out =  24'b000000000000000000011100;
		16'b1101100000110000 : data_out =  24'b000000000000000000011100;
		16'b1101100000110010 : data_out =  24'b000000000000000000011100;
		16'b1101100000110100 : data_out =  24'b000000000000000000011100;
		16'b1101100000110110 : data_out =  24'b000000000000000000011100;
		16'b1101100000111000 : data_out =  24'b000000000000000000011100;
		16'b1101100000111010 : data_out =  24'b000000000000000000011100;
		16'b1101100000111100 : data_out =  24'b000000000000000000011100;
		16'b1101100000111110 : data_out =  24'b000000000000000000011100;
		16'b1101100001000000 : data_out =  24'b000000000000000000011100;
		16'b1101100001000010 : data_out =  24'b000000000000000000011100;
		16'b1101100001000100 : data_out =  24'b000000000000000000011100;
		16'b1101100001000110 : data_out =  24'b000000000000000000011100;
		16'b1101100001001000 : data_out =  24'b000000000000000000011100;
		16'b1101100001001010 : data_out =  24'b000000000000000000011100;
		16'b1101100001001100 : data_out =  24'b000000000000000000011100;
		16'b1101100001001110 : data_out =  24'b000000000000000000011100;
		16'b1101100001010000 : data_out =  24'b000000000000000000011100;
		16'b1101100001010010 : data_out =  24'b000000000000000000011100;
		16'b1101100001010100 : data_out =  24'b000000000000000000011100;
		16'b1101100001010111 : data_out =  24'b000000000000000000011100;
		16'b1101100001011001 : data_out =  24'b000000000000000000011100;
		16'b1101100001011011 : data_out =  24'b000000000000000000011100;
		16'b1101100001011101 : data_out =  24'b000000000000000000011100;
		16'b1101100001011111 : data_out =  24'b000000000000000000011100;
		16'b1101100001100001 : data_out =  24'b000000000000000000011100;
		16'b1101100001100011 : data_out =  24'b000000000000000000011100;
		16'b1101100001100101 : data_out =  24'b000000000000000000011100;
		16'b1101100001100111 : data_out =  24'b000000000000000000011101;
		16'b1101100001101001 : data_out =  24'b000000000000000000011101;
		16'b1101100001101011 : data_out =  24'b000000000000000000011101;
		16'b1101100001101101 : data_out =  24'b000000000000000000011101;
		16'b1101100001101111 : data_out =  24'b000000000000000000011101;
		16'b1101100001110001 : data_out =  24'b000000000000000000011101;
		16'b1101100001110011 : data_out =  24'b000000000000000000011101;
		16'b1101100001110101 : data_out =  24'b000000000000000000011101;
		16'b1101100001110111 : data_out =  24'b000000000000000000011101;
		16'b1101100001111001 : data_out =  24'b000000000000000000011101;
		16'b1101100001111011 : data_out =  24'b000000000000000000011101;
		16'b1101100001111101 : data_out =  24'b000000000000000000011101;
		16'b1101100001111111 : data_out =  24'b000000000000000000011101;
		16'b1101100010000010 : data_out =  24'b000000000000000000011101;
		16'b1101100010000100 : data_out =  24'b000000000000000000011101;
		16'b1101100010000110 : data_out =  24'b000000000000000000011101;
		16'b1101100010001000 : data_out =  24'b000000000000000000011101;
		16'b1101100010001010 : data_out =  24'b000000000000000000011101;
		16'b1101100010001100 : data_out =  24'b000000000000000000011101;
		16'b1101100010001110 : data_out =  24'b000000000000000000011101;
		16'b1101100010010000 : data_out =  24'b000000000000000000011101;
		16'b1101100010010010 : data_out =  24'b000000000000000000011101;
		16'b1101100010010100 : data_out =  24'b000000000000000000011101;
		16'b1101100010010110 : data_out =  24'b000000000000000000011101;
		16'b1101100010011000 : data_out =  24'b000000000000000000011101;
		16'b1101100010011010 : data_out =  24'b000000000000000000011101;
		16'b1101100010011100 : data_out =  24'b000000000000000000011101;
		16'b1101100010011110 : data_out =  24'b000000000000000000011101;
		16'b1101100010100000 : data_out =  24'b000000000000000000011101;
		16'b1101100010100010 : data_out =  24'b000000000000000000011101;
		16'b1101100010100100 : data_out =  24'b000000000000000000011101;
		16'b1101100010100110 : data_out =  24'b000000000000000000011101;
		16'b1101100010101000 : data_out =  24'b000000000000000000011101;
		16'b1101100010101010 : data_out =  24'b000000000000000000011101;
		16'b1101100010101101 : data_out =  24'b000000000000000000011110;
		16'b1101100010101111 : data_out =  24'b000000000000000000011110;
		16'b1101100010110001 : data_out =  24'b000000000000000000011110;
		16'b1101100010110011 : data_out =  24'b000000000000000000011110;
		16'b1101100010110101 : data_out =  24'b000000000000000000011110;
		16'b1101100010110111 : data_out =  24'b000000000000000000011110;
		16'b1101100010111001 : data_out =  24'b000000000000000000011110;
		16'b1101100010111011 : data_out =  24'b000000000000000000011110;
		16'b1101100010111101 : data_out =  24'b000000000000000000011110;
		16'b1101100010111111 : data_out =  24'b000000000000000000011110;
		16'b1101100011000001 : data_out =  24'b000000000000000000011110;
		16'b1101100011000011 : data_out =  24'b000000000000000000011110;
		16'b1101100011000101 : data_out =  24'b000000000000000000011110;
		16'b1101100011000111 : data_out =  24'b000000000000000000011110;
		16'b1101100011001001 : data_out =  24'b000000000000000000011110;
		16'b1101100011001011 : data_out =  24'b000000000000000000011110;
		16'b1101100011001101 : data_out =  24'b000000000000000000011110;
		16'b1101100011001111 : data_out =  24'b000000000000000000011110;
		16'b1101100011010001 : data_out =  24'b000000000000000000011110;
		16'b1101100011010011 : data_out =  24'b000000000000000000011110;
		16'b1101100011010101 : data_out =  24'b000000000000000000011110;
		16'b1101100011011000 : data_out =  24'b000000000000000000011110;
		16'b1101100011011010 : data_out =  24'b000000000000000000011110;
		16'b1101100011011100 : data_out =  24'b000000000000000000011110;
		16'b1101100011011110 : data_out =  24'b000000000000000000011110;
		16'b1101100011100000 : data_out =  24'b000000000000000000011110;
		16'b1101100011100010 : data_out =  24'b000000000000000000011110;
		16'b1101100011100100 : data_out =  24'b000000000000000000011110;
		16'b1101100011100110 : data_out =  24'b000000000000000000011110;
		16'b1101100011101000 : data_out =  24'b000000000000000000011110;
		16'b1101100011101010 : data_out =  24'b000000000000000000011110;
		16'b1101100011101100 : data_out =  24'b000000000000000000011110;
		16'b1101100011101110 : data_out =  24'b000000000000000000011110;
		16'b1101100011110000 : data_out =  24'b000000000000000000011111;
		16'b1101100011110010 : data_out =  24'b000000000000000000011111;
		16'b1101100011110100 : data_out =  24'b000000000000000000011111;
		16'b1101100011110110 : data_out =  24'b000000000000000000011111;
		16'b1101100011111000 : data_out =  24'b000000000000000000011111;
		16'b1101100011111010 : data_out =  24'b000000000000000000011111;
		16'b1101100011111100 : data_out =  24'b000000000000000000011111;
		16'b1101100011111110 : data_out =  24'b000000000000000000011111;
		16'b1101100100000001 : data_out =  24'b000000000000000000011111;
		16'b1101100100000011 : data_out =  24'b000000000000000000011111;
		16'b1101100100000101 : data_out =  24'b000000000000000000011111;
		16'b1101100100000111 : data_out =  24'b000000000000000000011111;
		16'b1101100100001001 : data_out =  24'b000000000000000000011111;
		16'b1101100100001011 : data_out =  24'b000000000000000000011111;
		16'b1101100100001101 : data_out =  24'b000000000000000000011111;
		16'b1101100100001111 : data_out =  24'b000000000000000000011111;
		16'b1101100100010001 : data_out =  24'b000000000000000000011111;
		16'b1101100100010011 : data_out =  24'b000000000000000000011111;
		16'b1101100100010101 : data_out =  24'b000000000000000000011111;
		16'b1101100100010111 : data_out =  24'b000000000000000000011111;
		16'b1101100100011001 : data_out =  24'b000000000000000000011111;
		16'b1101100100011011 : data_out =  24'b000000000000000000011111;
		16'b1101100100011101 : data_out =  24'b000000000000000000011111;
		16'b1101100100011111 : data_out =  24'b000000000000000000011111;
		16'b1101100100100001 : data_out =  24'b000000000000000000011111;
		16'b1101100100100011 : data_out =  24'b000000000000000000011111;
		16'b1101100100100101 : data_out =  24'b000000000000000000011111;
		16'b1101100100100111 : data_out =  24'b000000000000000000011111;
		16'b1101100100101001 : data_out =  24'b000000000000000000011111;
		16'b1101100100101100 : data_out =  24'b000000000000000000011111;
		16'b1101100100101110 : data_out =  24'b000000000000000000011111;
		16'b1101100100110000 : data_out =  24'b000000000000000000100000;
		16'b1101100100110010 : data_out =  24'b000000000000000000100000;
		16'b1101100100110100 : data_out =  24'b000000000000000000100000;
		16'b1101100100110110 : data_out =  24'b000000000000000000100000;
		16'b1101100100111000 : data_out =  24'b000000000000000000100000;
		16'b1101100100111010 : data_out =  24'b000000000000000000100000;
		16'b1101100100111100 : data_out =  24'b000000000000000000100000;
		16'b1101100100111110 : data_out =  24'b000000000000000000100000;
		16'b1101100101000000 : data_out =  24'b000000000000000000100000;
		16'b1101100101000010 : data_out =  24'b000000000000000000100000;
		16'b1101100101000100 : data_out =  24'b000000000000000000100000;
		16'b1101100101000110 : data_out =  24'b000000000000000000100000;
		16'b1101100101001000 : data_out =  24'b000000000000000000100000;
		16'b1101100101001010 : data_out =  24'b000000000000000000100000;
		16'b1101100101001100 : data_out =  24'b000000000000000000100000;
		16'b1101100101001110 : data_out =  24'b000000000000000000100000;
		16'b1101100101010000 : data_out =  24'b000000000000000000100000;
		16'b1101100101010010 : data_out =  24'b000000000000000000100000;
		16'b1101100101010100 : data_out =  24'b000000000000000000100000;
		16'b1101100101010111 : data_out =  24'b000000000000000000100000;
		16'b1101100101011001 : data_out =  24'b000000000000000000100000;
		16'b1101100101011011 : data_out =  24'b000000000000000000100000;
		16'b1101100101011101 : data_out =  24'b000000000000000000100000;
		16'b1101100101011111 : data_out =  24'b000000000000000000100000;
		16'b1101100101100001 : data_out =  24'b000000000000000000100000;
		16'b1101100101100011 : data_out =  24'b000000000000000000100000;
		16'b1101100101100101 : data_out =  24'b000000000000000000100000;
		16'b1101100101100111 : data_out =  24'b000000000000000000100000;
		16'b1101100101101001 : data_out =  24'b000000000000000000100000;
		16'b1101100101101011 : data_out =  24'b000000000000000000100000;
		16'b1101100101101101 : data_out =  24'b000000000000000000100000;
		16'b1101100101101111 : data_out =  24'b000000000000000000100001;
		16'b1101100101110001 : data_out =  24'b000000000000000000100001;
		16'b1101100101110011 : data_out =  24'b000000000000000000100001;
		16'b1101100101110101 : data_out =  24'b000000000000000000100001;
		16'b1101100101110111 : data_out =  24'b000000000000000000100001;
		16'b1101100101111001 : data_out =  24'b000000000000000000100001;
		16'b1101100101111011 : data_out =  24'b000000000000000000100001;
		16'b1101100101111101 : data_out =  24'b000000000000000000100001;
		16'b1101100101111111 : data_out =  24'b000000000000000000100001;
		16'b1101100110000010 : data_out =  24'b000000000000000000100001;
		16'b1101100110000100 : data_out =  24'b000000000000000000100001;
		16'b1101100110000110 : data_out =  24'b000000000000000000100001;
		16'b1101100110001000 : data_out =  24'b000000000000000000100001;
		16'b1101100110001010 : data_out =  24'b000000000000000000100001;
		16'b1101100110001100 : data_out =  24'b000000000000000000100001;
		16'b1101100110001110 : data_out =  24'b000000000000000000100001;
		16'b1101100110010000 : data_out =  24'b000000000000000000100001;
		16'b1101100110010010 : data_out =  24'b000000000000000000100001;
		16'b1101100110010100 : data_out =  24'b000000000000000000100001;
		16'b1101100110010110 : data_out =  24'b000000000000000000100001;
		16'b1101100110011000 : data_out =  24'b000000000000000000100001;
		16'b1101100110011010 : data_out =  24'b000000000000000000100001;
		16'b1101100110011100 : data_out =  24'b000000000000000000100001;
		16'b1101100110011110 : data_out =  24'b000000000000000000100001;
		16'b1101100110100000 : data_out =  24'b000000000000000000100001;
		16'b1101100110100010 : data_out =  24'b000000000000000000100001;
		16'b1101100110100100 : data_out =  24'b000000000000000000100001;
		16'b1101100110100110 : data_out =  24'b000000000000000000100001;
		16'b1101100110101000 : data_out =  24'b000000000000000000100001;
		16'b1101100110101010 : data_out =  24'b000000000000000000100001;
		16'b1101100110101101 : data_out =  24'b000000000000000000100010;
		16'b1101100110101111 : data_out =  24'b000000000000000000100010;
		16'b1101100110110001 : data_out =  24'b000000000000000000100010;
		16'b1101100110110011 : data_out =  24'b000000000000000000100010;
		16'b1101100110110101 : data_out =  24'b000000000000000000100010;
		16'b1101100110110111 : data_out =  24'b000000000000000000100010;
		16'b1101100110111001 : data_out =  24'b000000000000000000100010;
		16'b1101100110111011 : data_out =  24'b000000000000000000100010;
		16'b1101100110111101 : data_out =  24'b000000000000000000100010;
		16'b1101100110111111 : data_out =  24'b000000000000000000100010;
		16'b1101100111000001 : data_out =  24'b000000000000000000100010;
		16'b1101100111000011 : data_out =  24'b000000000000000000100010;
		16'b1101100111000101 : data_out =  24'b000000000000000000100010;
		16'b1101100111000111 : data_out =  24'b000000000000000000100010;
		16'b1101100111001001 : data_out =  24'b000000000000000000100010;
		16'b1101100111001011 : data_out =  24'b000000000000000000100010;
		16'b1101100111001101 : data_out =  24'b000000000000000000100010;
		16'b1101100111001111 : data_out =  24'b000000000000000000100010;
		16'b1101100111010001 : data_out =  24'b000000000000000000100010;
		16'b1101100111010011 : data_out =  24'b000000000000000000100010;
		16'b1101100111010101 : data_out =  24'b000000000000000000100010;
		16'b1101100111011000 : data_out =  24'b000000000000000000100010;
		16'b1101100111011010 : data_out =  24'b000000000000000000100010;
		16'b1101100111011100 : data_out =  24'b000000000000000000100010;
		16'b1101100111011110 : data_out =  24'b000000000000000000100010;
		16'b1101100111100000 : data_out =  24'b000000000000000000100010;
		16'b1101100111100010 : data_out =  24'b000000000000000000100010;
		16'b1101100111100100 : data_out =  24'b000000000000000000100010;
		16'b1101100111100110 : data_out =  24'b000000000000000000100010;
		16'b1101100111101000 : data_out =  24'b000000000000000000100011;
		16'b1101100111101010 : data_out =  24'b000000000000000000100011;
		16'b1101100111101100 : data_out =  24'b000000000000000000100011;
		16'b1101100111101110 : data_out =  24'b000000000000000000100011;
		16'b1101100111110000 : data_out =  24'b000000000000000000100011;
		16'b1101100111110010 : data_out =  24'b000000000000000000100011;
		16'b1101100111110100 : data_out =  24'b000000000000000000100011;
		16'b1101100111110110 : data_out =  24'b000000000000000000100011;
		16'b1101100111111000 : data_out =  24'b000000000000000000100011;
		16'b1101100111111010 : data_out =  24'b000000000000000000100011;
		16'b1101100111111100 : data_out =  24'b000000000000000000100011;
		16'b1101100111111110 : data_out =  24'b000000000000000000100011;
		16'b1101101000000001 : data_out =  24'b000000000000000000100011;
		16'b1101101000000011 : data_out =  24'b000000000000000000100011;
		16'b1101101000000101 : data_out =  24'b000000000000000000100011;
		16'b1101101000000111 : data_out =  24'b000000000000000000100011;
		16'b1101101000001001 : data_out =  24'b000000000000000000100011;
		16'b1101101000001011 : data_out =  24'b000000000000000000100011;
		16'b1101101000001101 : data_out =  24'b000000000000000000100011;
		16'b1101101000001111 : data_out =  24'b000000000000000000100011;
		16'b1101101000010001 : data_out =  24'b000000000000000000100011;
		16'b1101101000010011 : data_out =  24'b000000000000000000100011;
		16'b1101101000010101 : data_out =  24'b000000000000000000100011;
		16'b1101101000010111 : data_out =  24'b000000000000000000100011;
		16'b1101101000011001 : data_out =  24'b000000000000000000100011;
		16'b1101101000011011 : data_out =  24'b000000000000000000100011;
		16'b1101101000011101 : data_out =  24'b000000000000000000100011;
		16'b1101101000011111 : data_out =  24'b000000000000000000100011;
		16'b1101101000100001 : data_out =  24'b000000000000000000100100;
		16'b1101101000100011 : data_out =  24'b000000000000000000100100;
		16'b1101101000100101 : data_out =  24'b000000000000000000100100;
		16'b1101101000100111 : data_out =  24'b000000000000000000100100;
		16'b1101101000101001 : data_out =  24'b000000000000000000100100;
		16'b1101101000101100 : data_out =  24'b000000000000000000100100;
		16'b1101101000101110 : data_out =  24'b000000000000000000100100;
		16'b1101101000110000 : data_out =  24'b000000000000000000100100;
		16'b1101101000110010 : data_out =  24'b000000000000000000100100;
		16'b1101101000110100 : data_out =  24'b000000000000000000100100;
		16'b1101101000110110 : data_out =  24'b000000000000000000100100;
		16'b1101101000111000 : data_out =  24'b000000000000000000100100;
		16'b1101101000111010 : data_out =  24'b000000000000000000100100;
		16'b1101101000111100 : data_out =  24'b000000000000000000100100;
		16'b1101101000111110 : data_out =  24'b000000000000000000100100;
		16'b1101101001000000 : data_out =  24'b000000000000000000100100;
		16'b1101101001000010 : data_out =  24'b000000000000000000100100;
		16'b1101101001000100 : data_out =  24'b000000000000000000100100;
		16'b1101101001000110 : data_out =  24'b000000000000000000100100;
		16'b1101101001001000 : data_out =  24'b000000000000000000100100;
		16'b1101101001001010 : data_out =  24'b000000000000000000100100;
		16'b1101101001001100 : data_out =  24'b000000000000000000100100;
		16'b1101101001001110 : data_out =  24'b000000000000000000100100;
		16'b1101101001010000 : data_out =  24'b000000000000000000100100;
		16'b1101101001010010 : data_out =  24'b000000000000000000100100;
		16'b1101101001010100 : data_out =  24'b000000000000000000100100;
		16'b1101101001010111 : data_out =  24'b000000000000000000100100;
		16'b1101101001011001 : data_out =  24'b000000000000000000100100;
		16'b1101101001011011 : data_out =  24'b000000000000000000100101;
		16'b1101101001011101 : data_out =  24'b000000000000000000100101;
		16'b1101101001011111 : data_out =  24'b000000000000000000100101;
		16'b1101101001100001 : data_out =  24'b000000000000000000100101;
		16'b1101101001100011 : data_out =  24'b000000000000000000100101;
		16'b1101101001100101 : data_out =  24'b000000000000000000100101;
		16'b1101101001100111 : data_out =  24'b000000000000000000100101;
		16'b1101101001101001 : data_out =  24'b000000000000000000100101;
		16'b1101101001101011 : data_out =  24'b000000000000000000100101;
		16'b1101101001101101 : data_out =  24'b000000000000000000100101;
		16'b1101101001101111 : data_out =  24'b000000000000000000100101;
		16'b1101101001110001 : data_out =  24'b000000000000000000100101;
		16'b1101101001110011 : data_out =  24'b000000000000000000100101;
		16'b1101101001110101 : data_out =  24'b000000000000000000100101;
		16'b1101101001110111 : data_out =  24'b000000000000000000100101;
		16'b1101101001111001 : data_out =  24'b000000000000000000100101;
		16'b1101101001111011 : data_out =  24'b000000000000000000100101;
		16'b1101101001111101 : data_out =  24'b000000000000000000100101;
		16'b1101101001111111 : data_out =  24'b000000000000000000100101;
		16'b1101101010000010 : data_out =  24'b000000000000000000100101;
		16'b1101101010000100 : data_out =  24'b000000000000000000100101;
		16'b1101101010000110 : data_out =  24'b000000000000000000100101;
		16'b1101101010001000 : data_out =  24'b000000000000000000100101;
		16'b1101101010001010 : data_out =  24'b000000000000000000100101;
		16'b1101101010001100 : data_out =  24'b000000000000000000100101;
		16'b1101101010001110 : data_out =  24'b000000000000000000100101;
		16'b1101101010010000 : data_out =  24'b000000000000000000100110;
		16'b1101101010010010 : data_out =  24'b000000000000000000100110;
		16'b1101101010010100 : data_out =  24'b000000000000000000100110;
		16'b1101101010010110 : data_out =  24'b000000000000000000100110;
		16'b1101101010011000 : data_out =  24'b000000000000000000100110;
		16'b1101101010011010 : data_out =  24'b000000000000000000100110;
		16'b1101101010011100 : data_out =  24'b000000000000000000100110;
		16'b1101101010011110 : data_out =  24'b000000000000000000100110;
		16'b1101101010100000 : data_out =  24'b000000000000000000100110;
		16'b1101101010100010 : data_out =  24'b000000000000000000100110;
		16'b1101101010100100 : data_out =  24'b000000000000000000100110;
		16'b1101101010100110 : data_out =  24'b000000000000000000100110;
		16'b1101101010101000 : data_out =  24'b000000000000000000100110;
		16'b1101101010101010 : data_out =  24'b000000000000000000100110;
		16'b1101101010101101 : data_out =  24'b000000000000000000100110;
		16'b1101101010101111 : data_out =  24'b000000000000000000100110;
		16'b1101101010110001 : data_out =  24'b000000000000000000100110;
		16'b1101101010110011 : data_out =  24'b000000000000000000100110;
		16'b1101101010110101 : data_out =  24'b000000000000000000100110;
		16'b1101101010110111 : data_out =  24'b000000000000000000100110;
		16'b1101101010111001 : data_out =  24'b000000000000000000100110;
		16'b1101101010111011 : data_out =  24'b000000000000000000100110;
		16'b1101101010111101 : data_out =  24'b000000000000000000100110;
		16'b1101101010111111 : data_out =  24'b000000000000000000100110;
		16'b1101101011000001 : data_out =  24'b000000000000000000100110;
		16'b1101101011000011 : data_out =  24'b000000000000000000100110;
		16'b1101101011000101 : data_out =  24'b000000000000000000100111;
		16'b1101101011000111 : data_out =  24'b000000000000000000100111;
		16'b1101101011001001 : data_out =  24'b000000000000000000100111;
		16'b1101101011001011 : data_out =  24'b000000000000000000100111;
		16'b1101101011001101 : data_out =  24'b000000000000000000100111;
		16'b1101101011001111 : data_out =  24'b000000000000000000100111;
		16'b1101101011010001 : data_out =  24'b000000000000000000100111;
		16'b1101101011010011 : data_out =  24'b000000000000000000100111;
		16'b1101101011010101 : data_out =  24'b000000000000000000100111;
		16'b1101101011011000 : data_out =  24'b000000000000000000100111;
		16'b1101101011011010 : data_out =  24'b000000000000000000100111;
		16'b1101101011011100 : data_out =  24'b000000000000000000100111;
		16'b1101101011011110 : data_out =  24'b000000000000000000100111;
		16'b1101101011100000 : data_out =  24'b000000000000000000100111;
		16'b1101101011100010 : data_out =  24'b000000000000000000100111;
		16'b1101101011100100 : data_out =  24'b000000000000000000100111;
		16'b1101101011100110 : data_out =  24'b000000000000000000100111;
		16'b1101101011101000 : data_out =  24'b000000000000000000100111;
		16'b1101101011101010 : data_out =  24'b000000000000000000100111;
		16'b1101101011101100 : data_out =  24'b000000000000000000100111;
		16'b1101101011101110 : data_out =  24'b000000000000000000100111;
		16'b1101101011110000 : data_out =  24'b000000000000000000100111;
		16'b1101101011110010 : data_out =  24'b000000000000000000100111;
		16'b1101101011110100 : data_out =  24'b000000000000000000100111;
		16'b1101101011110110 : data_out =  24'b000000000000000000100111;
		16'b1101101011111000 : data_out =  24'b000000000000000000100111;
		16'b1101101011111010 : data_out =  24'b000000000000000000101000;
		16'b1101101011111100 : data_out =  24'b000000000000000000101000;
		16'b1101101011111110 : data_out =  24'b000000000000000000101000;
		16'b1101101100000001 : data_out =  24'b000000000000000000101000;
		16'b1101101100000011 : data_out =  24'b000000000000000000101000;
		16'b1101101100000101 : data_out =  24'b000000000000000000101000;
		16'b1101101100000111 : data_out =  24'b000000000000000000101000;
		16'b1101101100001001 : data_out =  24'b000000000000000000101000;
		16'b1101101100001011 : data_out =  24'b000000000000000000101000;
		16'b1101101100001101 : data_out =  24'b000000000000000000101000;
		16'b1101101100001111 : data_out =  24'b000000000000000000101000;
		16'b1101101100010001 : data_out =  24'b000000000000000000101000;
		16'b1101101100010011 : data_out =  24'b000000000000000000101000;
		16'b1101101100010101 : data_out =  24'b000000000000000000101000;
		16'b1101101100010111 : data_out =  24'b000000000000000000101000;
		16'b1101101100011001 : data_out =  24'b000000000000000000101000;
		16'b1101101100011011 : data_out =  24'b000000000000000000101000;
		16'b1101101100011101 : data_out =  24'b000000000000000000101000;
		16'b1101101100011111 : data_out =  24'b000000000000000000101000;
		16'b1101101100100001 : data_out =  24'b000000000000000000101000;
		16'b1101101100100011 : data_out =  24'b000000000000000000101000;
		16'b1101101100100101 : data_out =  24'b000000000000000000101000;
		16'b1101101100100111 : data_out =  24'b000000000000000000101000;
		16'b1101101100101001 : data_out =  24'b000000000000000000101000;
		16'b1101101100101100 : data_out =  24'b000000000000000000101001;
		16'b1101101100101110 : data_out =  24'b000000000000000000101001;
		16'b1101101100110000 : data_out =  24'b000000000000000000101001;
		16'b1101101100110010 : data_out =  24'b000000000000000000101001;
		16'b1101101100110100 : data_out =  24'b000000000000000000101001;
		16'b1101101100110110 : data_out =  24'b000000000000000000101001;
		16'b1101101100111000 : data_out =  24'b000000000000000000101001;
		16'b1101101100111010 : data_out =  24'b000000000000000000101001;
		16'b1101101100111100 : data_out =  24'b000000000000000000101001;
		16'b1101101100111110 : data_out =  24'b000000000000000000101001;
		16'b1101101101000000 : data_out =  24'b000000000000000000101001;
		16'b1101101101000010 : data_out =  24'b000000000000000000101001;
		16'b1101101101000100 : data_out =  24'b000000000000000000101001;
		16'b1101101101000110 : data_out =  24'b000000000000000000101001;
		16'b1101101101001000 : data_out =  24'b000000000000000000101001;
		16'b1101101101001010 : data_out =  24'b000000000000000000101001;
		16'b1101101101001100 : data_out =  24'b000000000000000000101001;
		16'b1101101101001110 : data_out =  24'b000000000000000000101001;
		16'b1101101101010000 : data_out =  24'b000000000000000000101001;
		16'b1101101101010010 : data_out =  24'b000000000000000000101001;
		16'b1101101101010100 : data_out =  24'b000000000000000000101001;
		16'b1101101101010111 : data_out =  24'b000000000000000000101001;
		16'b1101101101011001 : data_out =  24'b000000000000000000101001;
		16'b1101101101011011 : data_out =  24'b000000000000000000101001;
		16'b1101101101011101 : data_out =  24'b000000000000000000101010;
		16'b1101101101011111 : data_out =  24'b000000000000000000101010;
		16'b1101101101100001 : data_out =  24'b000000000000000000101010;
		16'b1101101101100011 : data_out =  24'b000000000000000000101010;
		16'b1101101101100101 : data_out =  24'b000000000000000000101010;
		16'b1101101101100111 : data_out =  24'b000000000000000000101010;
		16'b1101101101101001 : data_out =  24'b000000000000000000101010;
		16'b1101101101101011 : data_out =  24'b000000000000000000101010;
		16'b1101101101101101 : data_out =  24'b000000000000000000101010;
		16'b1101101101101111 : data_out =  24'b000000000000000000101010;
		16'b1101101101110001 : data_out =  24'b000000000000000000101010;
		16'b1101101101110011 : data_out =  24'b000000000000000000101010;
		16'b1101101101110101 : data_out =  24'b000000000000000000101010;
		16'b1101101101110111 : data_out =  24'b000000000000000000101010;
		16'b1101101101111001 : data_out =  24'b000000000000000000101010;
		16'b1101101101111011 : data_out =  24'b000000000000000000101010;
		16'b1101101101111101 : data_out =  24'b000000000000000000101010;
		16'b1101101101111111 : data_out =  24'b000000000000000000101010;
		16'b1101101110000010 : data_out =  24'b000000000000000000101010;
		16'b1101101110000100 : data_out =  24'b000000000000000000101010;
		16'b1101101110000110 : data_out =  24'b000000000000000000101010;
		16'b1101101110001000 : data_out =  24'b000000000000000000101010;
		16'b1101101110001010 : data_out =  24'b000000000000000000101010;
		16'b1101101110001100 : data_out =  24'b000000000000000000101010;
		16'b1101101110001110 : data_out =  24'b000000000000000000101011;
		16'b1101101110010000 : data_out =  24'b000000000000000000101011;
		16'b1101101110010010 : data_out =  24'b000000000000000000101011;
		16'b1101101110010100 : data_out =  24'b000000000000000000101011;
		16'b1101101110010110 : data_out =  24'b000000000000000000101011;
		16'b1101101110011000 : data_out =  24'b000000000000000000101011;
		16'b1101101110011010 : data_out =  24'b000000000000000000101011;
		16'b1101101110011100 : data_out =  24'b000000000000000000101011;
		16'b1101101110011110 : data_out =  24'b000000000000000000101011;
		16'b1101101110100000 : data_out =  24'b000000000000000000101011;
		16'b1101101110100010 : data_out =  24'b000000000000000000101011;
		16'b1101101110100100 : data_out =  24'b000000000000000000101011;
		16'b1101101110100110 : data_out =  24'b000000000000000000101011;
		16'b1101101110101000 : data_out =  24'b000000000000000000101011;
		16'b1101101110101010 : data_out =  24'b000000000000000000101011;
		16'b1101101110101101 : data_out =  24'b000000000000000000101011;
		16'b1101101110101111 : data_out =  24'b000000000000000000101011;
		16'b1101101110110001 : data_out =  24'b000000000000000000101011;
		16'b1101101110110011 : data_out =  24'b000000000000000000101011;
		16'b1101101110110101 : data_out =  24'b000000000000000000101011;
		16'b1101101110110111 : data_out =  24'b000000000000000000101011;
		16'b1101101110111001 : data_out =  24'b000000000000000000101011;
		16'b1101101110111011 : data_out =  24'b000000000000000000101011;
		16'b1101101110111101 : data_out =  24'b000000000000000000101100;
		16'b1101101110111111 : data_out =  24'b000000000000000000101100;
		16'b1101101111000001 : data_out =  24'b000000000000000000101100;
		16'b1101101111000011 : data_out =  24'b000000000000000000101100;
		16'b1101101111000101 : data_out =  24'b000000000000000000101100;
		16'b1101101111000111 : data_out =  24'b000000000000000000101100;
		16'b1101101111001001 : data_out =  24'b000000000000000000101100;
		16'b1101101111001011 : data_out =  24'b000000000000000000101100;
		16'b1101101111001101 : data_out =  24'b000000000000000000101100;
		16'b1101101111001111 : data_out =  24'b000000000000000000101100;
		16'b1101101111010001 : data_out =  24'b000000000000000000101100;
		16'b1101101111010011 : data_out =  24'b000000000000000000101100;
		16'b1101101111010101 : data_out =  24'b000000000000000000101100;
		16'b1101101111011000 : data_out =  24'b000000000000000000101100;
		16'b1101101111011010 : data_out =  24'b000000000000000000101100;
		16'b1101101111011100 : data_out =  24'b000000000000000000101100;
		16'b1101101111011110 : data_out =  24'b000000000000000000101100;
		16'b1101101111100000 : data_out =  24'b000000000000000000101100;
		16'b1101101111100010 : data_out =  24'b000000000000000000101100;
		16'b1101101111100100 : data_out =  24'b000000000000000000101100;
		16'b1101101111100110 : data_out =  24'b000000000000000000101100;
		16'b1101101111101000 : data_out =  24'b000000000000000000101100;
		16'b1101101111101010 : data_out =  24'b000000000000000000101101;
		16'b1101101111101100 : data_out =  24'b000000000000000000101101;
		16'b1101101111101110 : data_out =  24'b000000000000000000101101;
		16'b1101101111110000 : data_out =  24'b000000000000000000101101;
		16'b1101101111110010 : data_out =  24'b000000000000000000101101;
		16'b1101101111110100 : data_out =  24'b000000000000000000101101;
		16'b1101101111110110 : data_out =  24'b000000000000000000101101;
		16'b1101101111111000 : data_out =  24'b000000000000000000101101;
		16'b1101101111111010 : data_out =  24'b000000000000000000101101;
		16'b1101101111111100 : data_out =  24'b000000000000000000101101;
		16'b1101101111111110 : data_out =  24'b000000000000000000101101;
		16'b1101110000000001 : data_out =  24'b000000000000000000101101;
		16'b1101110000000011 : data_out =  24'b000000000000000000101101;
		16'b1101110000000101 : data_out =  24'b000000000000000000101101;
		16'b1101110000000111 : data_out =  24'b000000000000000000101101;
		16'b1101110000001001 : data_out =  24'b000000000000000000101101;
		16'b1101110000001011 : data_out =  24'b000000000000000000101101;
		16'b1101110000001101 : data_out =  24'b000000000000000000101101;
		16'b1101110000001111 : data_out =  24'b000000000000000000101101;
		16'b1101110000010001 : data_out =  24'b000000000000000000101101;
		16'b1101110000010011 : data_out =  24'b000000000000000000101101;
		16'b1101110000010101 : data_out =  24'b000000000000000000101101;
		16'b1101110000010111 : data_out =  24'b000000000000000000101110;
		16'b1101110000011001 : data_out =  24'b000000000000000000101110;
		16'b1101110000011011 : data_out =  24'b000000000000000000101110;
		16'b1101110000011101 : data_out =  24'b000000000000000000101110;
		16'b1101110000011111 : data_out =  24'b000000000000000000101110;
		16'b1101110000100001 : data_out =  24'b000000000000000000101110;
		16'b1101110000100011 : data_out =  24'b000000000000000000101110;
		16'b1101110000100101 : data_out =  24'b000000000000000000101110;
		16'b1101110000100111 : data_out =  24'b000000000000000000101110;
		16'b1101110000101001 : data_out =  24'b000000000000000000101110;
		16'b1101110000101100 : data_out =  24'b000000000000000000101110;
		16'b1101110000101110 : data_out =  24'b000000000000000000101110;
		16'b1101110000110000 : data_out =  24'b000000000000000000101110;
		16'b1101110000110010 : data_out =  24'b000000000000000000101110;
		16'b1101110000110100 : data_out =  24'b000000000000000000101110;
		16'b1101110000110110 : data_out =  24'b000000000000000000101110;
		16'b1101110000111000 : data_out =  24'b000000000000000000101110;
		16'b1101110000111010 : data_out =  24'b000000000000000000101110;
		16'b1101110000111100 : data_out =  24'b000000000000000000101110;
		16'b1101110000111110 : data_out =  24'b000000000000000000101110;
		16'b1101110001000000 : data_out =  24'b000000000000000000101110;
		16'b1101110001000010 : data_out =  24'b000000000000000000101110;
		16'b1101110001000100 : data_out =  24'b000000000000000000101111;
		16'b1101110001000110 : data_out =  24'b000000000000000000101111;
		16'b1101110001001000 : data_out =  24'b000000000000000000101111;
		16'b1101110001001010 : data_out =  24'b000000000000000000101111;
		16'b1101110001001100 : data_out =  24'b000000000000000000101111;
		16'b1101110001001110 : data_out =  24'b000000000000000000101111;
		16'b1101110001010000 : data_out =  24'b000000000000000000101111;
		16'b1101110001010010 : data_out =  24'b000000000000000000101111;
		16'b1101110001010100 : data_out =  24'b000000000000000000101111;
		16'b1101110001010111 : data_out =  24'b000000000000000000101111;
		16'b1101110001011001 : data_out =  24'b000000000000000000101111;
		16'b1101110001011011 : data_out =  24'b000000000000000000101111;
		16'b1101110001011101 : data_out =  24'b000000000000000000101111;
		16'b1101110001011111 : data_out =  24'b000000000000000000101111;
		16'b1101110001100001 : data_out =  24'b000000000000000000101111;
		16'b1101110001100011 : data_out =  24'b000000000000000000101111;
		16'b1101110001100101 : data_out =  24'b000000000000000000101111;
		16'b1101110001100111 : data_out =  24'b000000000000000000101111;
		16'b1101110001101001 : data_out =  24'b000000000000000000101111;
		16'b1101110001101011 : data_out =  24'b000000000000000000101111;
		16'b1101110001101101 : data_out =  24'b000000000000000000101111;
		16'b1101110001101111 : data_out =  24'b000000000000000000110000;
		16'b1101110001110001 : data_out =  24'b000000000000000000110000;
		16'b1101110001110011 : data_out =  24'b000000000000000000110000;
		16'b1101110001110101 : data_out =  24'b000000000000000000110000;
		16'b1101110001110111 : data_out =  24'b000000000000000000110000;
		16'b1101110001111001 : data_out =  24'b000000000000000000110000;
		16'b1101110001111011 : data_out =  24'b000000000000000000110000;
		16'b1101110001111101 : data_out =  24'b000000000000000000110000;
		16'b1101110001111111 : data_out =  24'b000000000000000000110000;
		16'b1101110010000010 : data_out =  24'b000000000000000000110000;
		16'b1101110010000100 : data_out =  24'b000000000000000000110000;
		16'b1101110010000110 : data_out =  24'b000000000000000000110000;
		16'b1101110010001000 : data_out =  24'b000000000000000000110000;
		16'b1101110010001010 : data_out =  24'b000000000000000000110000;
		16'b1101110010001100 : data_out =  24'b000000000000000000110000;
		16'b1101110010001110 : data_out =  24'b000000000000000000110000;
		16'b1101110010010000 : data_out =  24'b000000000000000000110000;
		16'b1101110010010010 : data_out =  24'b000000000000000000110000;
		16'b1101110010010100 : data_out =  24'b000000000000000000110000;
		16'b1101110010010110 : data_out =  24'b000000000000000000110000;
		16'b1101110010011000 : data_out =  24'b000000000000000000110000;
		16'b1101110010011010 : data_out =  24'b000000000000000000110001;
		16'b1101110010011100 : data_out =  24'b000000000000000000110001;
		16'b1101110010011110 : data_out =  24'b000000000000000000110001;
		16'b1101110010100000 : data_out =  24'b000000000000000000110001;
		16'b1101110010100010 : data_out =  24'b000000000000000000110001;
		16'b1101110010100100 : data_out =  24'b000000000000000000110001;
		16'b1101110010100110 : data_out =  24'b000000000000000000110001;
		16'b1101110010101000 : data_out =  24'b000000000000000000110001;
		16'b1101110010101010 : data_out =  24'b000000000000000000110001;
		16'b1101110010101101 : data_out =  24'b000000000000000000110001;
		16'b1101110010101111 : data_out =  24'b000000000000000000110001;
		16'b1101110010110001 : data_out =  24'b000000000000000000110001;
		16'b1101110010110011 : data_out =  24'b000000000000000000110001;
		16'b1101110010110101 : data_out =  24'b000000000000000000110001;
		16'b1101110010110111 : data_out =  24'b000000000000000000110001;
		16'b1101110010111001 : data_out =  24'b000000000000000000110001;
		16'b1101110010111011 : data_out =  24'b000000000000000000110001;
		16'b1101110010111101 : data_out =  24'b000000000000000000110001;
		16'b1101110010111111 : data_out =  24'b000000000000000000110001;
		16'b1101110011000001 : data_out =  24'b000000000000000000110001;
		16'b1101110011000011 : data_out =  24'b000000000000000000110010;
		16'b1101110011000101 : data_out =  24'b000000000000000000110010;
		16'b1101110011000111 : data_out =  24'b000000000000000000110010;
		16'b1101110011001001 : data_out =  24'b000000000000000000110010;
		16'b1101110011001011 : data_out =  24'b000000000000000000110010;
		16'b1101110011001101 : data_out =  24'b000000000000000000110010;
		16'b1101110011001111 : data_out =  24'b000000000000000000110010;
		16'b1101110011010001 : data_out =  24'b000000000000000000110010;
		16'b1101110011010011 : data_out =  24'b000000000000000000110010;
		16'b1101110011010101 : data_out =  24'b000000000000000000110010;
		16'b1101110011011000 : data_out =  24'b000000000000000000110010;
		16'b1101110011011010 : data_out =  24'b000000000000000000110010;
		16'b1101110011011100 : data_out =  24'b000000000000000000110010;
		16'b1101110011011110 : data_out =  24'b000000000000000000110010;
		16'b1101110011100000 : data_out =  24'b000000000000000000110010;
		16'b1101110011100010 : data_out =  24'b000000000000000000110010;
		16'b1101110011100100 : data_out =  24'b000000000000000000110010;
		16'b1101110011100110 : data_out =  24'b000000000000000000110010;
		16'b1101110011101000 : data_out =  24'b000000000000000000110010;
		16'b1101110011101010 : data_out =  24'b000000000000000000110010;
		16'b1101110011101100 : data_out =  24'b000000000000000000110011;
		16'b1101110011101110 : data_out =  24'b000000000000000000110011;
		16'b1101110011110000 : data_out =  24'b000000000000000000110011;
		16'b1101110011110010 : data_out =  24'b000000000000000000110011;
		16'b1101110011110100 : data_out =  24'b000000000000000000110011;
		16'b1101110011110110 : data_out =  24'b000000000000000000110011;
		16'b1101110011111000 : data_out =  24'b000000000000000000110011;
		16'b1101110011111010 : data_out =  24'b000000000000000000110011;
		16'b1101110011111100 : data_out =  24'b000000000000000000110011;
		16'b1101110011111110 : data_out =  24'b000000000000000000110011;
		16'b1101110100000001 : data_out =  24'b000000000000000000110011;
		16'b1101110100000011 : data_out =  24'b000000000000000000110011;
		16'b1101110100000101 : data_out =  24'b000000000000000000110011;
		16'b1101110100000111 : data_out =  24'b000000000000000000110011;
		16'b1101110100001001 : data_out =  24'b000000000000000000110011;
		16'b1101110100001011 : data_out =  24'b000000000000000000110011;
		16'b1101110100001101 : data_out =  24'b000000000000000000110011;
		16'b1101110100001111 : data_out =  24'b000000000000000000110011;
		16'b1101110100010001 : data_out =  24'b000000000000000000110011;
		16'b1101110100010011 : data_out =  24'b000000000000000000110100;
		16'b1101110100010101 : data_out =  24'b000000000000000000110100;
		16'b1101110100010111 : data_out =  24'b000000000000000000110100;
		16'b1101110100011001 : data_out =  24'b000000000000000000110100;
		16'b1101110100011011 : data_out =  24'b000000000000000000110100;
		16'b1101110100011101 : data_out =  24'b000000000000000000110100;
		16'b1101110100011111 : data_out =  24'b000000000000000000110100;
		16'b1101110100100001 : data_out =  24'b000000000000000000110100;
		16'b1101110100100011 : data_out =  24'b000000000000000000110100;
		16'b1101110100100101 : data_out =  24'b000000000000000000110100;
		16'b1101110100100111 : data_out =  24'b000000000000000000110100;
		16'b1101110100101001 : data_out =  24'b000000000000000000110100;
		16'b1101110100101100 : data_out =  24'b000000000000000000110100;
		16'b1101110100101110 : data_out =  24'b000000000000000000110100;
		16'b1101110100110000 : data_out =  24'b000000000000000000110100;
		16'b1101110100110010 : data_out =  24'b000000000000000000110100;
		16'b1101110100110100 : data_out =  24'b000000000000000000110100;
		16'b1101110100110110 : data_out =  24'b000000000000000000110100;
		16'b1101110100111000 : data_out =  24'b000000000000000000110100;
		16'b1101110100111010 : data_out =  24'b000000000000000000110101;
		16'b1101110100111100 : data_out =  24'b000000000000000000110101;
		16'b1101110100111110 : data_out =  24'b000000000000000000110101;
		16'b1101110101000000 : data_out =  24'b000000000000000000110101;
		16'b1101110101000010 : data_out =  24'b000000000000000000110101;
		16'b1101110101000100 : data_out =  24'b000000000000000000110101;
		16'b1101110101000110 : data_out =  24'b000000000000000000110101;
		16'b1101110101001000 : data_out =  24'b000000000000000000110101;
		16'b1101110101001010 : data_out =  24'b000000000000000000110101;
		16'b1101110101001100 : data_out =  24'b000000000000000000110101;
		16'b1101110101001110 : data_out =  24'b000000000000000000110101;
		16'b1101110101010000 : data_out =  24'b000000000000000000110101;
		16'b1101110101010010 : data_out =  24'b000000000000000000110101;
		16'b1101110101010100 : data_out =  24'b000000000000000000110101;
		16'b1101110101010111 : data_out =  24'b000000000000000000110101;
		16'b1101110101011001 : data_out =  24'b000000000000000000110101;
		16'b1101110101011011 : data_out =  24'b000000000000000000110101;
		16'b1101110101011101 : data_out =  24'b000000000000000000110101;
		16'b1101110101011111 : data_out =  24'b000000000000000000110101;
		16'b1101110101100001 : data_out =  24'b000000000000000000110110;
		16'b1101110101100011 : data_out =  24'b000000000000000000110110;
		16'b1101110101100101 : data_out =  24'b000000000000000000110110;
		16'b1101110101100111 : data_out =  24'b000000000000000000110110;
		16'b1101110101101001 : data_out =  24'b000000000000000000110110;
		16'b1101110101101011 : data_out =  24'b000000000000000000110110;
		16'b1101110101101101 : data_out =  24'b000000000000000000110110;
		16'b1101110101101111 : data_out =  24'b000000000000000000110110;
		16'b1101110101110001 : data_out =  24'b000000000000000000110110;
		16'b1101110101110011 : data_out =  24'b000000000000000000110110;
		16'b1101110101110101 : data_out =  24'b000000000000000000110110;
		16'b1101110101110111 : data_out =  24'b000000000000000000110110;
		16'b1101110101111001 : data_out =  24'b000000000000000000110110;
		16'b1101110101111011 : data_out =  24'b000000000000000000110110;
		16'b1101110101111101 : data_out =  24'b000000000000000000110110;
		16'b1101110101111111 : data_out =  24'b000000000000000000110110;
		16'b1101110110000010 : data_out =  24'b000000000000000000110110;
		16'b1101110110000100 : data_out =  24'b000000000000000000110110;
		16'b1101110110000110 : data_out =  24'b000000000000000000110111;
		16'b1101110110001000 : data_out =  24'b000000000000000000110111;
		16'b1101110110001010 : data_out =  24'b000000000000000000110111;
		16'b1101110110001100 : data_out =  24'b000000000000000000110111;
		16'b1101110110001110 : data_out =  24'b000000000000000000110111;
		16'b1101110110010000 : data_out =  24'b000000000000000000110111;
		16'b1101110110010010 : data_out =  24'b000000000000000000110111;
		16'b1101110110010100 : data_out =  24'b000000000000000000110111;
		16'b1101110110010110 : data_out =  24'b000000000000000000110111;
		16'b1101110110011000 : data_out =  24'b000000000000000000110111;
		16'b1101110110011010 : data_out =  24'b000000000000000000110111;
		16'b1101110110011100 : data_out =  24'b000000000000000000110111;
		16'b1101110110011110 : data_out =  24'b000000000000000000110111;
		16'b1101110110100000 : data_out =  24'b000000000000000000110111;
		16'b1101110110100010 : data_out =  24'b000000000000000000110111;
		16'b1101110110100100 : data_out =  24'b000000000000000000110111;
		16'b1101110110100110 : data_out =  24'b000000000000000000110111;
		16'b1101110110101000 : data_out =  24'b000000000000000000110111;
		16'b1101110110101010 : data_out =  24'b000000000000000000111000;
		16'b1101110110101101 : data_out =  24'b000000000000000000111000;
		16'b1101110110101111 : data_out =  24'b000000000000000000111000;
		16'b1101110110110001 : data_out =  24'b000000000000000000111000;
		16'b1101110110110011 : data_out =  24'b000000000000000000111000;
		16'b1101110110110101 : data_out =  24'b000000000000000000111000;
		16'b1101110110110111 : data_out =  24'b000000000000000000111000;
		16'b1101110110111001 : data_out =  24'b000000000000000000111000;
		16'b1101110110111011 : data_out =  24'b000000000000000000111000;
		16'b1101110110111101 : data_out =  24'b000000000000000000111000;
		16'b1101110110111111 : data_out =  24'b000000000000000000111000;
		16'b1101110111000001 : data_out =  24'b000000000000000000111000;
		16'b1101110111000011 : data_out =  24'b000000000000000000111000;
		16'b1101110111000101 : data_out =  24'b000000000000000000111000;
		16'b1101110111000111 : data_out =  24'b000000000000000000111000;
		16'b1101110111001001 : data_out =  24'b000000000000000000111000;
		16'b1101110111001011 : data_out =  24'b000000000000000000111000;
		16'b1101110111001101 : data_out =  24'b000000000000000000111000;
		16'b1101110111001111 : data_out =  24'b000000000000000000111001;
		16'b1101110111010001 : data_out =  24'b000000000000000000111001;
		16'b1101110111010011 : data_out =  24'b000000000000000000111001;
		16'b1101110111010101 : data_out =  24'b000000000000000000111001;
		16'b1101110111011000 : data_out =  24'b000000000000000000111001;
		16'b1101110111011010 : data_out =  24'b000000000000000000111001;
		16'b1101110111011100 : data_out =  24'b000000000000000000111001;
		16'b1101110111011110 : data_out =  24'b000000000000000000111001;
		16'b1101110111100000 : data_out =  24'b000000000000000000111001;
		16'b1101110111100010 : data_out =  24'b000000000000000000111001;
		16'b1101110111100100 : data_out =  24'b000000000000000000111001;
		16'b1101110111100110 : data_out =  24'b000000000000000000111001;
		16'b1101110111101000 : data_out =  24'b000000000000000000111001;
		16'b1101110111101010 : data_out =  24'b000000000000000000111001;
		16'b1101110111101100 : data_out =  24'b000000000000000000111001;
		16'b1101110111101110 : data_out =  24'b000000000000000000111001;
		16'b1101110111110000 : data_out =  24'b000000000000000000111001;
		16'b1101110111110010 : data_out =  24'b000000000000000000111010;
		16'b1101110111110100 : data_out =  24'b000000000000000000111010;
		16'b1101110111110110 : data_out =  24'b000000000000000000111010;
		16'b1101110111111000 : data_out =  24'b000000000000000000111010;
		16'b1101110111111010 : data_out =  24'b000000000000000000111010;
		16'b1101110111111100 : data_out =  24'b000000000000000000111010;
		16'b1101110111111110 : data_out =  24'b000000000000000000111010;
		16'b1101111000000001 : data_out =  24'b000000000000000000111010;
		16'b1101111000000011 : data_out =  24'b000000000000000000111010;
		16'b1101111000000101 : data_out =  24'b000000000000000000111010;
		16'b1101111000000111 : data_out =  24'b000000000000000000111010;
		16'b1101111000001001 : data_out =  24'b000000000000000000111010;
		16'b1101111000001011 : data_out =  24'b000000000000000000111010;
		16'b1101111000001101 : data_out =  24'b000000000000000000111010;
		16'b1101111000001111 : data_out =  24'b000000000000000000111010;
		16'b1101111000010001 : data_out =  24'b000000000000000000111010;
		16'b1101111000010011 : data_out =  24'b000000000000000000111010;
		16'b1101111000010101 : data_out =  24'b000000000000000000111011;
		16'b1101111000010111 : data_out =  24'b000000000000000000111011;
		16'b1101111000011001 : data_out =  24'b000000000000000000111011;
		16'b1101111000011011 : data_out =  24'b000000000000000000111011;
		16'b1101111000011101 : data_out =  24'b000000000000000000111011;
		16'b1101111000011111 : data_out =  24'b000000000000000000111011;
		16'b1101111000100001 : data_out =  24'b000000000000000000111011;
		16'b1101111000100011 : data_out =  24'b000000000000000000111011;
		16'b1101111000100101 : data_out =  24'b000000000000000000111011;
		16'b1101111000100111 : data_out =  24'b000000000000000000111011;
		16'b1101111000101001 : data_out =  24'b000000000000000000111011;
		16'b1101111000101100 : data_out =  24'b000000000000000000111011;
		16'b1101111000101110 : data_out =  24'b000000000000000000111011;
		16'b1101111000110000 : data_out =  24'b000000000000000000111011;
		16'b1101111000110010 : data_out =  24'b000000000000000000111011;
		16'b1101111000110100 : data_out =  24'b000000000000000000111011;
		16'b1101111000110110 : data_out =  24'b000000000000000000111011;
		16'b1101111000111000 : data_out =  24'b000000000000000000111100;
		16'b1101111000111010 : data_out =  24'b000000000000000000111100;
		16'b1101111000111100 : data_out =  24'b000000000000000000111100;
		16'b1101111000111110 : data_out =  24'b000000000000000000111100;
		16'b1101111001000000 : data_out =  24'b000000000000000000111100;
		16'b1101111001000010 : data_out =  24'b000000000000000000111100;
		16'b1101111001000100 : data_out =  24'b000000000000000000111100;
		16'b1101111001000110 : data_out =  24'b000000000000000000111100;
		16'b1101111001001000 : data_out =  24'b000000000000000000111100;
		16'b1101111001001010 : data_out =  24'b000000000000000000111100;
		16'b1101111001001100 : data_out =  24'b000000000000000000111100;
		16'b1101111001001110 : data_out =  24'b000000000000000000111100;
		16'b1101111001010000 : data_out =  24'b000000000000000000111100;
		16'b1101111001010010 : data_out =  24'b000000000000000000111100;
		16'b1101111001010100 : data_out =  24'b000000000000000000111100;
		16'b1101111001010111 : data_out =  24'b000000000000000000111100;
		16'b1101111001011001 : data_out =  24'b000000000000000000111100;
		16'b1101111001011011 : data_out =  24'b000000000000000000111101;
		16'b1101111001011101 : data_out =  24'b000000000000000000111101;
		16'b1101111001011111 : data_out =  24'b000000000000000000111101;
		16'b1101111001100001 : data_out =  24'b000000000000000000111101;
		16'b1101111001100011 : data_out =  24'b000000000000000000111101;
		16'b1101111001100101 : data_out =  24'b000000000000000000111101;
		16'b1101111001100111 : data_out =  24'b000000000000000000111101;
		16'b1101111001101001 : data_out =  24'b000000000000000000111101;
		16'b1101111001101011 : data_out =  24'b000000000000000000111101;
		16'b1101111001101101 : data_out =  24'b000000000000000000111101;
		16'b1101111001101111 : data_out =  24'b000000000000000000111101;
		16'b1101111001110001 : data_out =  24'b000000000000000000111101;
		16'b1101111001110011 : data_out =  24'b000000000000000000111101;
		16'b1101111001110101 : data_out =  24'b000000000000000000111101;
		16'b1101111001110111 : data_out =  24'b000000000000000000111101;
		16'b1101111001111001 : data_out =  24'b000000000000000000111101;
		16'b1101111001111011 : data_out =  24'b000000000000000000111110;
		16'b1101111001111101 : data_out =  24'b000000000000000000111110;
		16'b1101111001111111 : data_out =  24'b000000000000000000111110;
		16'b1101111010000010 : data_out =  24'b000000000000000000111110;
		16'b1101111010000100 : data_out =  24'b000000000000000000111110;
		16'b1101111010000110 : data_out =  24'b000000000000000000111110;
		16'b1101111010001000 : data_out =  24'b000000000000000000111110;
		16'b1101111010001010 : data_out =  24'b000000000000000000111110;
		16'b1101111010001100 : data_out =  24'b000000000000000000111110;
		16'b1101111010001110 : data_out =  24'b000000000000000000111110;
		16'b1101111010010000 : data_out =  24'b000000000000000000111110;
		16'b1101111010010010 : data_out =  24'b000000000000000000111110;
		16'b1101111010010100 : data_out =  24'b000000000000000000111110;
		16'b1101111010010110 : data_out =  24'b000000000000000000111110;
		16'b1101111010011000 : data_out =  24'b000000000000000000111110;
		16'b1101111010011010 : data_out =  24'b000000000000000000111110;
		16'b1101111010011100 : data_out =  24'b000000000000000000111111;
		16'b1101111010011110 : data_out =  24'b000000000000000000111111;
		16'b1101111010100000 : data_out =  24'b000000000000000000111111;
		16'b1101111010100010 : data_out =  24'b000000000000000000111111;
		16'b1101111010100100 : data_out =  24'b000000000000000000111111;
		16'b1101111010100110 : data_out =  24'b000000000000000000111111;
		16'b1101111010101000 : data_out =  24'b000000000000000000111111;
		16'b1101111010101010 : data_out =  24'b000000000000000000111111;
		16'b1101111010101101 : data_out =  24'b000000000000000000111111;
		16'b1101111010101111 : data_out =  24'b000000000000000000111111;
		16'b1101111010110001 : data_out =  24'b000000000000000000111111;
		16'b1101111010110011 : data_out =  24'b000000000000000000111111;
		16'b1101111010110101 : data_out =  24'b000000000000000000111111;
		16'b1101111010110111 : data_out =  24'b000000000000000000111111;
		16'b1101111010111001 : data_out =  24'b000000000000000000111111;
		16'b1101111010111011 : data_out =  24'b000000000000000000111111;
		16'b1101111010111101 : data_out =  24'b000000000000000001000000;
		16'b1101111010111111 : data_out =  24'b000000000000000001000000;
		16'b1101111011000001 : data_out =  24'b000000000000000001000000;
		16'b1101111011000011 : data_out =  24'b000000000000000001000000;
		16'b1101111011000101 : data_out =  24'b000000000000000001000000;
		16'b1101111011000111 : data_out =  24'b000000000000000001000000;
		16'b1101111011001001 : data_out =  24'b000000000000000001000000;
		16'b1101111011001011 : data_out =  24'b000000000000000001000000;
		16'b1101111011001101 : data_out =  24'b000000000000000001000000;
		16'b1101111011001111 : data_out =  24'b000000000000000001000000;
		16'b1101111011010001 : data_out =  24'b000000000000000001000000;
		16'b1101111011010011 : data_out =  24'b000000000000000001000000;
		16'b1101111011010101 : data_out =  24'b000000000000000001000000;
		16'b1101111011011000 : data_out =  24'b000000000000000001000000;
		16'b1101111011011010 : data_out =  24'b000000000000000001000000;
		16'b1101111011011100 : data_out =  24'b000000000000000001000001;
		16'b1101111011011110 : data_out =  24'b000000000000000001000001;
		16'b1101111011100000 : data_out =  24'b000000000000000001000001;
		16'b1101111011100010 : data_out =  24'b000000000000000001000001;
		16'b1101111011100100 : data_out =  24'b000000000000000001000001;
		16'b1101111011100110 : data_out =  24'b000000000000000001000001;
		16'b1101111011101000 : data_out =  24'b000000000000000001000001;
		16'b1101111011101010 : data_out =  24'b000000000000000001000001;
		16'b1101111011101100 : data_out =  24'b000000000000000001000001;
		16'b1101111011101110 : data_out =  24'b000000000000000001000001;
		16'b1101111011110000 : data_out =  24'b000000000000000001000001;
		16'b1101111011110010 : data_out =  24'b000000000000000001000001;
		16'b1101111011110100 : data_out =  24'b000000000000000001000001;
		16'b1101111011110110 : data_out =  24'b000000000000000001000001;
		16'b1101111011111000 : data_out =  24'b000000000000000001000001;
		16'b1101111011111010 : data_out =  24'b000000000000000001000010;
		16'b1101111011111100 : data_out =  24'b000000000000000001000010;
		16'b1101111011111110 : data_out =  24'b000000000000000001000010;
		16'b1101111100000001 : data_out =  24'b000000000000000001000010;
		16'b1101111100000011 : data_out =  24'b000000000000000001000010;
		16'b1101111100000101 : data_out =  24'b000000000000000001000010;
		16'b1101111100000111 : data_out =  24'b000000000000000001000010;
		16'b1101111100001001 : data_out =  24'b000000000000000001000010;
		16'b1101111100001011 : data_out =  24'b000000000000000001000010;
		16'b1101111100001101 : data_out =  24'b000000000000000001000010;
		16'b1101111100001111 : data_out =  24'b000000000000000001000010;
		16'b1101111100010001 : data_out =  24'b000000000000000001000010;
		16'b1101111100010011 : data_out =  24'b000000000000000001000010;
		16'b1101111100010101 : data_out =  24'b000000000000000001000010;
		16'b1101111100010111 : data_out =  24'b000000000000000001000010;
		16'b1101111100011001 : data_out =  24'b000000000000000001000011;
		16'b1101111100011011 : data_out =  24'b000000000000000001000011;
		16'b1101111100011101 : data_out =  24'b000000000000000001000011;
		16'b1101111100011111 : data_out =  24'b000000000000000001000011;
		16'b1101111100100001 : data_out =  24'b000000000000000001000011;
		16'b1101111100100011 : data_out =  24'b000000000000000001000011;
		16'b1101111100100101 : data_out =  24'b000000000000000001000011;
		16'b1101111100100111 : data_out =  24'b000000000000000001000011;
		16'b1101111100101001 : data_out =  24'b000000000000000001000011;
		16'b1101111100101100 : data_out =  24'b000000000000000001000011;
		16'b1101111100101110 : data_out =  24'b000000000000000001000011;
		16'b1101111100110000 : data_out =  24'b000000000000000001000011;
		16'b1101111100110010 : data_out =  24'b000000000000000001000011;
		16'b1101111100110100 : data_out =  24'b000000000000000001000011;
		16'b1101111100110110 : data_out =  24'b000000000000000001000011;
		16'b1101111100111000 : data_out =  24'b000000000000000001000100;
		16'b1101111100111010 : data_out =  24'b000000000000000001000100;
		16'b1101111100111100 : data_out =  24'b000000000000000001000100;
		16'b1101111100111110 : data_out =  24'b000000000000000001000100;
		16'b1101111101000000 : data_out =  24'b000000000000000001000100;
		16'b1101111101000010 : data_out =  24'b000000000000000001000100;
		16'b1101111101000100 : data_out =  24'b000000000000000001000100;
		16'b1101111101000110 : data_out =  24'b000000000000000001000100;
		16'b1101111101001000 : data_out =  24'b000000000000000001000100;
		16'b1101111101001010 : data_out =  24'b000000000000000001000100;
		16'b1101111101001100 : data_out =  24'b000000000000000001000100;
		16'b1101111101001110 : data_out =  24'b000000000000000001000100;
		16'b1101111101010000 : data_out =  24'b000000000000000001000100;
		16'b1101111101010010 : data_out =  24'b000000000000000001000100;
		16'b1101111101010100 : data_out =  24'b000000000000000001000100;
		16'b1101111101010111 : data_out =  24'b000000000000000001000101;
		16'b1101111101011001 : data_out =  24'b000000000000000001000101;
		16'b1101111101011011 : data_out =  24'b000000000000000001000101;
		16'b1101111101011101 : data_out =  24'b000000000000000001000101;
		16'b1101111101011111 : data_out =  24'b000000000000000001000101;
		16'b1101111101100001 : data_out =  24'b000000000000000001000101;
		16'b1101111101100011 : data_out =  24'b000000000000000001000101;
		16'b1101111101100101 : data_out =  24'b000000000000000001000101;
		16'b1101111101100111 : data_out =  24'b000000000000000001000101;
		16'b1101111101101001 : data_out =  24'b000000000000000001000101;
		16'b1101111101101011 : data_out =  24'b000000000000000001000101;
		16'b1101111101101101 : data_out =  24'b000000000000000001000101;
		16'b1101111101101111 : data_out =  24'b000000000000000001000101;
		16'b1101111101110001 : data_out =  24'b000000000000000001000101;
		16'b1101111101110011 : data_out =  24'b000000000000000001000110;
		16'b1101111101110101 : data_out =  24'b000000000000000001000110;
		16'b1101111101110111 : data_out =  24'b000000000000000001000110;
		16'b1101111101111001 : data_out =  24'b000000000000000001000110;
		16'b1101111101111011 : data_out =  24'b000000000000000001000110;
		16'b1101111101111101 : data_out =  24'b000000000000000001000110;
		16'b1101111101111111 : data_out =  24'b000000000000000001000110;
		16'b1101111110000010 : data_out =  24'b000000000000000001000110;
		16'b1101111110000100 : data_out =  24'b000000000000000001000110;
		16'b1101111110000110 : data_out =  24'b000000000000000001000110;
		16'b1101111110001000 : data_out =  24'b000000000000000001000110;
		16'b1101111110001010 : data_out =  24'b000000000000000001000110;
		16'b1101111110001100 : data_out =  24'b000000000000000001000110;
		16'b1101111110001110 : data_out =  24'b000000000000000001000110;
		16'b1101111110010000 : data_out =  24'b000000000000000001000111;
		16'b1101111110010010 : data_out =  24'b000000000000000001000111;
		16'b1101111110010100 : data_out =  24'b000000000000000001000111;
		16'b1101111110010110 : data_out =  24'b000000000000000001000111;
		16'b1101111110011000 : data_out =  24'b000000000000000001000111;
		16'b1101111110011010 : data_out =  24'b000000000000000001000111;
		16'b1101111110011100 : data_out =  24'b000000000000000001000111;
		16'b1101111110011110 : data_out =  24'b000000000000000001000111;
		16'b1101111110100000 : data_out =  24'b000000000000000001000111;
		16'b1101111110100010 : data_out =  24'b000000000000000001000111;
		16'b1101111110100100 : data_out =  24'b000000000000000001000111;
		16'b1101111110100110 : data_out =  24'b000000000000000001000111;
		16'b1101111110101000 : data_out =  24'b000000000000000001000111;
		16'b1101111110101010 : data_out =  24'b000000000000000001000111;
		16'b1101111110101101 : data_out =  24'b000000000000000001001000;
		16'b1101111110101111 : data_out =  24'b000000000000000001001000;
		16'b1101111110110001 : data_out =  24'b000000000000000001001000;
		16'b1101111110110011 : data_out =  24'b000000000000000001001000;
		16'b1101111110110101 : data_out =  24'b000000000000000001001000;
		16'b1101111110110111 : data_out =  24'b000000000000000001001000;
		16'b1101111110111001 : data_out =  24'b000000000000000001001000;
		16'b1101111110111011 : data_out =  24'b000000000000000001001000;
		16'b1101111110111101 : data_out =  24'b000000000000000001001000;
		16'b1101111110111111 : data_out =  24'b000000000000000001001000;
		16'b1101111111000001 : data_out =  24'b000000000000000001001000;
		16'b1101111111000011 : data_out =  24'b000000000000000001001000;
		16'b1101111111000101 : data_out =  24'b000000000000000001001000;
		16'b1101111111000111 : data_out =  24'b000000000000000001001000;
		16'b1101111111001001 : data_out =  24'b000000000000000001001001;
		16'b1101111111001011 : data_out =  24'b000000000000000001001001;
		16'b1101111111001101 : data_out =  24'b000000000000000001001001;
		16'b1101111111001111 : data_out =  24'b000000000000000001001001;
		16'b1101111111010001 : data_out =  24'b000000000000000001001001;
		16'b1101111111010011 : data_out =  24'b000000000000000001001001;
		16'b1101111111010101 : data_out =  24'b000000000000000001001001;
		16'b1101111111011000 : data_out =  24'b000000000000000001001001;
		16'b1101111111011010 : data_out =  24'b000000000000000001001001;
		16'b1101111111011100 : data_out =  24'b000000000000000001001001;
		16'b1101111111011110 : data_out =  24'b000000000000000001001001;
		16'b1101111111100000 : data_out =  24'b000000000000000001001001;
		16'b1101111111100010 : data_out =  24'b000000000000000001001001;
		16'b1101111111100100 : data_out =  24'b000000000000000001001001;
		16'b1101111111100110 : data_out =  24'b000000000000000001001010;
		16'b1101111111101000 : data_out =  24'b000000000000000001001010;
		16'b1101111111101010 : data_out =  24'b000000000000000001001010;
		16'b1101111111101100 : data_out =  24'b000000000000000001001010;
		16'b1101111111101110 : data_out =  24'b000000000000000001001010;
		16'b1101111111110000 : data_out =  24'b000000000000000001001010;
		16'b1101111111110010 : data_out =  24'b000000000000000001001010;
		16'b1101111111110100 : data_out =  24'b000000000000000001001010;
		16'b1101111111110110 : data_out =  24'b000000000000000001001010;
		16'b1101111111111000 : data_out =  24'b000000000000000001001010;
		16'b1101111111111010 : data_out =  24'b000000000000000001001010;
		16'b1101111111111100 : data_out =  24'b000000000000000001001010;
		16'b1101111111111110 : data_out =  24'b000000000000000001001010;
		16'b1110000000000001 : data_out =  24'b000000000000000001001011;
		16'b1110000000000011 : data_out =  24'b000000000000000001001011;
		16'b1110000000000101 : data_out =  24'b000000000000000001001011;
		16'b1110000000000111 : data_out =  24'b000000000000000001001011;
		16'b1110000000001001 : data_out =  24'b000000000000000001001011;
		16'b1110000000001011 : data_out =  24'b000000000000000001001011;
		16'b1110000000001101 : data_out =  24'b000000000000000001001011;
		16'b1110000000001111 : data_out =  24'b000000000000000001001011;
		16'b1110000000010001 : data_out =  24'b000000000000000001001011;
		16'b1110000000010011 : data_out =  24'b000000000000000001001011;
		16'b1110000000010101 : data_out =  24'b000000000000000001001011;
		16'b1110000000010111 : data_out =  24'b000000000000000001001011;
		16'b1110000000011001 : data_out =  24'b000000000000000001001011;
		16'b1110000000011011 : data_out =  24'b000000000000000001001100;
		16'b1110000000011101 : data_out =  24'b000000000000000001001100;
		16'b1110000000011111 : data_out =  24'b000000000000000001001100;
		16'b1110000000100001 : data_out =  24'b000000000000000001001100;
		16'b1110000000100011 : data_out =  24'b000000000000000001001100;
		16'b1110000000100101 : data_out =  24'b000000000000000001001100;
		16'b1110000000100111 : data_out =  24'b000000000000000001001100;
		16'b1110000000101001 : data_out =  24'b000000000000000001001100;
		16'b1110000000101100 : data_out =  24'b000000000000000001001100;
		16'b1110000000101110 : data_out =  24'b000000000000000001001100;
		16'b1110000000110000 : data_out =  24'b000000000000000001001100;
		16'b1110000000110010 : data_out =  24'b000000000000000001001100;
		16'b1110000000110100 : data_out =  24'b000000000000000001001100;
		16'b1110000000110110 : data_out =  24'b000000000000000001001100;
		16'b1110000000111000 : data_out =  24'b000000000000000001001101;
		16'b1110000000111010 : data_out =  24'b000000000000000001001101;
		16'b1110000000111100 : data_out =  24'b000000000000000001001101;
		16'b1110000000111110 : data_out =  24'b000000000000000001001101;
		16'b1110000001000000 : data_out =  24'b000000000000000001001101;
		16'b1110000001000010 : data_out =  24'b000000000000000001001101;
		16'b1110000001000100 : data_out =  24'b000000000000000001001101;
		16'b1110000001000110 : data_out =  24'b000000000000000001001101;
		16'b1110000001001000 : data_out =  24'b000000000000000001001101;
		16'b1110000001001010 : data_out =  24'b000000000000000001001101;
		16'b1110000001001100 : data_out =  24'b000000000000000001001101;
		16'b1110000001001110 : data_out =  24'b000000000000000001001101;
		16'b1110000001010000 : data_out =  24'b000000000000000001001110;
		16'b1110000001010010 : data_out =  24'b000000000000000001001110;
		16'b1110000001010100 : data_out =  24'b000000000000000001001110;
		16'b1110000001010111 : data_out =  24'b000000000000000001001110;
		16'b1110000001011001 : data_out =  24'b000000000000000001001110;
		16'b1110000001011011 : data_out =  24'b000000000000000001001110;
		16'b1110000001011101 : data_out =  24'b000000000000000001001110;
		16'b1110000001011111 : data_out =  24'b000000000000000001001110;
		16'b1110000001100001 : data_out =  24'b000000000000000001001110;
		16'b1110000001100011 : data_out =  24'b000000000000000001001110;
		16'b1110000001100101 : data_out =  24'b000000000000000001001110;
		16'b1110000001100111 : data_out =  24'b000000000000000001001110;
		16'b1110000001101001 : data_out =  24'b000000000000000001001110;
		16'b1110000001101011 : data_out =  24'b000000000000000001001111;
		16'b1110000001101101 : data_out =  24'b000000000000000001001111;
		16'b1110000001101111 : data_out =  24'b000000000000000001001111;
		16'b1110000001110001 : data_out =  24'b000000000000000001001111;
		16'b1110000001110011 : data_out =  24'b000000000000000001001111;
		16'b1110000001110101 : data_out =  24'b000000000000000001001111;
		16'b1110000001110111 : data_out =  24'b000000000000000001001111;
		16'b1110000001111001 : data_out =  24'b000000000000000001001111;
		16'b1110000001111011 : data_out =  24'b000000000000000001001111;
		16'b1110000001111101 : data_out =  24'b000000000000000001001111;
		16'b1110000001111111 : data_out =  24'b000000000000000001001111;
		16'b1110000010000010 : data_out =  24'b000000000000000001001111;
		16'b1110000010000100 : data_out =  24'b000000000000000001001111;
		16'b1110000010000110 : data_out =  24'b000000000000000001010000;
		16'b1110000010001000 : data_out =  24'b000000000000000001010000;
		16'b1110000010001010 : data_out =  24'b000000000000000001010000;
		16'b1110000010001100 : data_out =  24'b000000000000000001010000;
		16'b1110000010001110 : data_out =  24'b000000000000000001010000;
		16'b1110000010010000 : data_out =  24'b000000000000000001010000;
		16'b1110000010010010 : data_out =  24'b000000000000000001010000;
		16'b1110000010010100 : data_out =  24'b000000000000000001010000;
		16'b1110000010010110 : data_out =  24'b000000000000000001010000;
		16'b1110000010011000 : data_out =  24'b000000000000000001010000;
		16'b1110000010011010 : data_out =  24'b000000000000000001010000;
		16'b1110000010011100 : data_out =  24'b000000000000000001010000;
		16'b1110000010011110 : data_out =  24'b000000000000000001010001;
		16'b1110000010100000 : data_out =  24'b000000000000000001010001;
		16'b1110000010100010 : data_out =  24'b000000000000000001010001;
		16'b1110000010100100 : data_out =  24'b000000000000000001010001;
		16'b1110000010100110 : data_out =  24'b000000000000000001010001;
		16'b1110000010101000 : data_out =  24'b000000000000000001010001;
		16'b1110000010101010 : data_out =  24'b000000000000000001010001;
		16'b1110000010101101 : data_out =  24'b000000000000000001010001;
		16'b1110000010101111 : data_out =  24'b000000000000000001010001;
		16'b1110000010110001 : data_out =  24'b000000000000000001010001;
		16'b1110000010110011 : data_out =  24'b000000000000000001010001;
		16'b1110000010110101 : data_out =  24'b000000000000000001010001;
		16'b1110000010110111 : data_out =  24'b000000000000000001010010;
		16'b1110000010111001 : data_out =  24'b000000000000000001010010;
		16'b1110000010111011 : data_out =  24'b000000000000000001010010;
		16'b1110000010111101 : data_out =  24'b000000000000000001010010;
		16'b1110000010111111 : data_out =  24'b000000000000000001010010;
		16'b1110000011000001 : data_out =  24'b000000000000000001010010;
		16'b1110000011000011 : data_out =  24'b000000000000000001010010;
		16'b1110000011000101 : data_out =  24'b000000000000000001010010;
		16'b1110000011000111 : data_out =  24'b000000000000000001010010;
		16'b1110000011001001 : data_out =  24'b000000000000000001010010;
		16'b1110000011001011 : data_out =  24'b000000000000000001010010;
		16'b1110000011001101 : data_out =  24'b000000000000000001010010;
		16'b1110000011001111 : data_out =  24'b000000000000000001010010;
		16'b1110000011010001 : data_out =  24'b000000000000000001010011;
		16'b1110000011010011 : data_out =  24'b000000000000000001010011;
		16'b1110000011010101 : data_out =  24'b000000000000000001010011;
		16'b1110000011011000 : data_out =  24'b000000000000000001010011;
		16'b1110000011011010 : data_out =  24'b000000000000000001010011;
		16'b1110000011011100 : data_out =  24'b000000000000000001010011;
		16'b1110000011011110 : data_out =  24'b000000000000000001010011;
		16'b1110000011100000 : data_out =  24'b000000000000000001010011;
		16'b1110000011100010 : data_out =  24'b000000000000000001010011;
		16'b1110000011100100 : data_out =  24'b000000000000000001010011;
		16'b1110000011100110 : data_out =  24'b000000000000000001010011;
		16'b1110000011101000 : data_out =  24'b000000000000000001010011;
		16'b1110000011101010 : data_out =  24'b000000000000000001010100;
		16'b1110000011101100 : data_out =  24'b000000000000000001010100;
		16'b1110000011101110 : data_out =  24'b000000000000000001010100;
		16'b1110000011110000 : data_out =  24'b000000000000000001010100;
		16'b1110000011110010 : data_out =  24'b000000000000000001010100;
		16'b1110000011110100 : data_out =  24'b000000000000000001010100;
		16'b1110000011110110 : data_out =  24'b000000000000000001010100;
		16'b1110000011111000 : data_out =  24'b000000000000000001010100;
		16'b1110000011111010 : data_out =  24'b000000000000000001010100;
		16'b1110000011111100 : data_out =  24'b000000000000000001010100;
		16'b1110000011111110 : data_out =  24'b000000000000000001010100;
		16'b1110000100000001 : data_out =  24'b000000000000000001010101;
		16'b1110000100000011 : data_out =  24'b000000000000000001010101;
		16'b1110000100000101 : data_out =  24'b000000000000000001010101;
		16'b1110000100000111 : data_out =  24'b000000000000000001010101;
		16'b1110000100001001 : data_out =  24'b000000000000000001010101;
		16'b1110000100001011 : data_out =  24'b000000000000000001010101;
		16'b1110000100001101 : data_out =  24'b000000000000000001010101;
		16'b1110000100001111 : data_out =  24'b000000000000000001010101;
		16'b1110000100010001 : data_out =  24'b000000000000000001010101;
		16'b1110000100010011 : data_out =  24'b000000000000000001010101;
		16'b1110000100010101 : data_out =  24'b000000000000000001010101;
		16'b1110000100010111 : data_out =  24'b000000000000000001010101;
		16'b1110000100011001 : data_out =  24'b000000000000000001010110;
		16'b1110000100011011 : data_out =  24'b000000000000000001010110;
		16'b1110000100011101 : data_out =  24'b000000000000000001010110;
		16'b1110000100011111 : data_out =  24'b000000000000000001010110;
		16'b1110000100100001 : data_out =  24'b000000000000000001010110;
		16'b1110000100100011 : data_out =  24'b000000000000000001010110;
		16'b1110000100100101 : data_out =  24'b000000000000000001010110;
		16'b1110000100100111 : data_out =  24'b000000000000000001010110;
		16'b1110000100101001 : data_out =  24'b000000000000000001010110;
		16'b1110000100101100 : data_out =  24'b000000000000000001010110;
		16'b1110000100101110 : data_out =  24'b000000000000000001010110;
		16'b1110000100110000 : data_out =  24'b000000000000000001010110;
		16'b1110000100110010 : data_out =  24'b000000000000000001010111;
		16'b1110000100110100 : data_out =  24'b000000000000000001010111;
		16'b1110000100110110 : data_out =  24'b000000000000000001010111;
		16'b1110000100111000 : data_out =  24'b000000000000000001010111;
		16'b1110000100111010 : data_out =  24'b000000000000000001010111;
		16'b1110000100111100 : data_out =  24'b000000000000000001010111;
		16'b1110000100111110 : data_out =  24'b000000000000000001010111;
		16'b1110000101000000 : data_out =  24'b000000000000000001010111;
		16'b1110000101000010 : data_out =  24'b000000000000000001010111;
		16'b1110000101000100 : data_out =  24'b000000000000000001010111;
		16'b1110000101000110 : data_out =  24'b000000000000000001010111;
		16'b1110000101001000 : data_out =  24'b000000000000000001011000;
		16'b1110000101001010 : data_out =  24'b000000000000000001011000;
		16'b1110000101001100 : data_out =  24'b000000000000000001011000;
		16'b1110000101001110 : data_out =  24'b000000000000000001011000;
		16'b1110000101010000 : data_out =  24'b000000000000000001011000;
		16'b1110000101010010 : data_out =  24'b000000000000000001011000;
		16'b1110000101010100 : data_out =  24'b000000000000000001011000;
		16'b1110000101010111 : data_out =  24'b000000000000000001011000;
		16'b1110000101011001 : data_out =  24'b000000000000000001011000;
		16'b1110000101011011 : data_out =  24'b000000000000000001011000;
		16'b1110000101011101 : data_out =  24'b000000000000000001011000;
		16'b1110000101011111 : data_out =  24'b000000000000000001011001;
		16'b1110000101100001 : data_out =  24'b000000000000000001011001;
		16'b1110000101100011 : data_out =  24'b000000000000000001011001;
		16'b1110000101100101 : data_out =  24'b000000000000000001011001;
		16'b1110000101100111 : data_out =  24'b000000000000000001011001;
		16'b1110000101101001 : data_out =  24'b000000000000000001011001;
		16'b1110000101101011 : data_out =  24'b000000000000000001011001;
		16'b1110000101101101 : data_out =  24'b000000000000000001011001;
		16'b1110000101101111 : data_out =  24'b000000000000000001011001;
		16'b1110000101110001 : data_out =  24'b000000000000000001011001;
		16'b1110000101110011 : data_out =  24'b000000000000000001011001;
		16'b1110000101110101 : data_out =  24'b000000000000000001011001;
		16'b1110000101110111 : data_out =  24'b000000000000000001011010;
		16'b1110000101111001 : data_out =  24'b000000000000000001011010;
		16'b1110000101111011 : data_out =  24'b000000000000000001011010;
		16'b1110000101111101 : data_out =  24'b000000000000000001011010;
		16'b1110000101111111 : data_out =  24'b000000000000000001011010;
		16'b1110000110000010 : data_out =  24'b000000000000000001011010;
		16'b1110000110000100 : data_out =  24'b000000000000000001011010;
		16'b1110000110000110 : data_out =  24'b000000000000000001011010;
		16'b1110000110001000 : data_out =  24'b000000000000000001011010;
		16'b1110000110001010 : data_out =  24'b000000000000000001011010;
		16'b1110000110001100 : data_out =  24'b000000000000000001011010;
		16'b1110000110001110 : data_out =  24'b000000000000000001011011;
		16'b1110000110010000 : data_out =  24'b000000000000000001011011;
		16'b1110000110010010 : data_out =  24'b000000000000000001011011;
		16'b1110000110010100 : data_out =  24'b000000000000000001011011;
		16'b1110000110010110 : data_out =  24'b000000000000000001011011;
		16'b1110000110011000 : data_out =  24'b000000000000000001011011;
		16'b1110000110011010 : data_out =  24'b000000000000000001011011;
		16'b1110000110011100 : data_out =  24'b000000000000000001011011;
		16'b1110000110011110 : data_out =  24'b000000000000000001011011;
		16'b1110000110100000 : data_out =  24'b000000000000000001011011;
		16'b1110000110100010 : data_out =  24'b000000000000000001011011;
		16'b1110000110100100 : data_out =  24'b000000000000000001011100;
		16'b1110000110100110 : data_out =  24'b000000000000000001011100;
		16'b1110000110101000 : data_out =  24'b000000000000000001011100;
		16'b1110000110101010 : data_out =  24'b000000000000000001011100;
		16'b1110000110101101 : data_out =  24'b000000000000000001011100;
		16'b1110000110101111 : data_out =  24'b000000000000000001011100;
		16'b1110000110110001 : data_out =  24'b000000000000000001011100;
		16'b1110000110110011 : data_out =  24'b000000000000000001011100;
		16'b1110000110110101 : data_out =  24'b000000000000000001011100;
		16'b1110000110110111 : data_out =  24'b000000000000000001011100;
		16'b1110000110111001 : data_out =  24'b000000000000000001011101;
		16'b1110000110111011 : data_out =  24'b000000000000000001011101;
		16'b1110000110111101 : data_out =  24'b000000000000000001011101;
		16'b1110000110111111 : data_out =  24'b000000000000000001011101;
		16'b1110000111000001 : data_out =  24'b000000000000000001011101;
		16'b1110000111000011 : data_out =  24'b000000000000000001011101;
		16'b1110000111000101 : data_out =  24'b000000000000000001011101;
		16'b1110000111000111 : data_out =  24'b000000000000000001011101;
		16'b1110000111001001 : data_out =  24'b000000000000000001011101;
		16'b1110000111001011 : data_out =  24'b000000000000000001011101;
		16'b1110000111001101 : data_out =  24'b000000000000000001011101;
		16'b1110000111001111 : data_out =  24'b000000000000000001011110;
		16'b1110000111010001 : data_out =  24'b000000000000000001011110;
		16'b1110000111010011 : data_out =  24'b000000000000000001011110;
		16'b1110000111010101 : data_out =  24'b000000000000000001011110;
		16'b1110000111011000 : data_out =  24'b000000000000000001011110;
		16'b1110000111011010 : data_out =  24'b000000000000000001011110;
		16'b1110000111011100 : data_out =  24'b000000000000000001011110;
		16'b1110000111011110 : data_out =  24'b000000000000000001011110;
		16'b1110000111100000 : data_out =  24'b000000000000000001011110;
		16'b1110000111100010 : data_out =  24'b000000000000000001011110;
		16'b1110000111100100 : data_out =  24'b000000000000000001011110;
		16'b1110000111100110 : data_out =  24'b000000000000000001011111;
		16'b1110000111101000 : data_out =  24'b000000000000000001011111;
		16'b1110000111101010 : data_out =  24'b000000000000000001011111;
		16'b1110000111101100 : data_out =  24'b000000000000000001011111;
		16'b1110000111101110 : data_out =  24'b000000000000000001011111;
		16'b1110000111110000 : data_out =  24'b000000000000000001011111;
		16'b1110000111110010 : data_out =  24'b000000000000000001011111;
		16'b1110000111110100 : data_out =  24'b000000000000000001011111;
		16'b1110000111110110 : data_out =  24'b000000000000000001011111;
		16'b1110000111111000 : data_out =  24'b000000000000000001011111;
		16'b1110000111111010 : data_out =  24'b000000000000000001100000;
		16'b1110000111111100 : data_out =  24'b000000000000000001100000;
		16'b1110000111111110 : data_out =  24'b000000000000000001100000;
		16'b1110001000000001 : data_out =  24'b000000000000000001100000;
		16'b1110001000000011 : data_out =  24'b000000000000000001100000;
		16'b1110001000000101 : data_out =  24'b000000000000000001100000;
		16'b1110001000000111 : data_out =  24'b000000000000000001100000;
		16'b1110001000001001 : data_out =  24'b000000000000000001100000;
		16'b1110001000001011 : data_out =  24'b000000000000000001100000;
		16'b1110001000001101 : data_out =  24'b000000000000000001100000;
		16'b1110001000001111 : data_out =  24'b000000000000000001100001;
		16'b1110001000010001 : data_out =  24'b000000000000000001100001;
		16'b1110001000010011 : data_out =  24'b000000000000000001100001;
		16'b1110001000010101 : data_out =  24'b000000000000000001100001;
		16'b1110001000010111 : data_out =  24'b000000000000000001100001;
		16'b1110001000011001 : data_out =  24'b000000000000000001100001;
		16'b1110001000011011 : data_out =  24'b000000000000000001100001;
		16'b1110001000011101 : data_out =  24'b000000000000000001100001;
		16'b1110001000011111 : data_out =  24'b000000000000000001100001;
		16'b1110001000100001 : data_out =  24'b000000000000000001100001;
		16'b1110001000100011 : data_out =  24'b000000000000000001100001;
		16'b1110001000100101 : data_out =  24'b000000000000000001100010;
		16'b1110001000100111 : data_out =  24'b000000000000000001100010;
		16'b1110001000101001 : data_out =  24'b000000000000000001100010;
		16'b1110001000101100 : data_out =  24'b000000000000000001100010;
		16'b1110001000101110 : data_out =  24'b000000000000000001100010;
		16'b1110001000110000 : data_out =  24'b000000000000000001100010;
		16'b1110001000110010 : data_out =  24'b000000000000000001100010;
		16'b1110001000110100 : data_out =  24'b000000000000000001100010;
		16'b1110001000110110 : data_out =  24'b000000000000000001100010;
		16'b1110001000111000 : data_out =  24'b000000000000000001100010;
		16'b1110001000111010 : data_out =  24'b000000000000000001100011;
		16'b1110001000111100 : data_out =  24'b000000000000000001100011;
		16'b1110001000111110 : data_out =  24'b000000000000000001100011;
		16'b1110001001000000 : data_out =  24'b000000000000000001100011;
		16'b1110001001000010 : data_out =  24'b000000000000000001100011;
		16'b1110001001000100 : data_out =  24'b000000000000000001100011;
		16'b1110001001000110 : data_out =  24'b000000000000000001100011;
		16'b1110001001001000 : data_out =  24'b000000000000000001100011;
		16'b1110001001001010 : data_out =  24'b000000000000000001100011;
		16'b1110001001001100 : data_out =  24'b000000000000000001100011;
		16'b1110001001001110 : data_out =  24'b000000000000000001100100;
		16'b1110001001010000 : data_out =  24'b000000000000000001100100;
		16'b1110001001010010 : data_out =  24'b000000000000000001100100;
		16'b1110001001010100 : data_out =  24'b000000000000000001100100;
		16'b1110001001010111 : data_out =  24'b000000000000000001100100;
		16'b1110001001011001 : data_out =  24'b000000000000000001100100;
		16'b1110001001011011 : data_out =  24'b000000000000000001100100;
		16'b1110001001011101 : data_out =  24'b000000000000000001100100;
		16'b1110001001011111 : data_out =  24'b000000000000000001100100;
		16'b1110001001100001 : data_out =  24'b000000000000000001100100;
		16'b1110001001100011 : data_out =  24'b000000000000000001100101;
		16'b1110001001100101 : data_out =  24'b000000000000000001100101;
		16'b1110001001100111 : data_out =  24'b000000000000000001100101;
		16'b1110001001101001 : data_out =  24'b000000000000000001100101;
		16'b1110001001101011 : data_out =  24'b000000000000000001100101;
		16'b1110001001101101 : data_out =  24'b000000000000000001100101;
		16'b1110001001101111 : data_out =  24'b000000000000000001100101;
		16'b1110001001110001 : data_out =  24'b000000000000000001100101;
		16'b1110001001110011 : data_out =  24'b000000000000000001100101;
		16'b1110001001110101 : data_out =  24'b000000000000000001100101;
		16'b1110001001110111 : data_out =  24'b000000000000000001100110;
		16'b1110001001111001 : data_out =  24'b000000000000000001100110;
		16'b1110001001111011 : data_out =  24'b000000000000000001100110;
		16'b1110001001111101 : data_out =  24'b000000000000000001100110;
		16'b1110001001111111 : data_out =  24'b000000000000000001100110;
		16'b1110001010000010 : data_out =  24'b000000000000000001100110;
		16'b1110001010000100 : data_out =  24'b000000000000000001100110;
		16'b1110001010000110 : data_out =  24'b000000000000000001100110;
		16'b1110001010001000 : data_out =  24'b000000000000000001100110;
		16'b1110001010001010 : data_out =  24'b000000000000000001100111;
		16'b1110001010001100 : data_out =  24'b000000000000000001100111;
		16'b1110001010001110 : data_out =  24'b000000000000000001100111;
		16'b1110001010010000 : data_out =  24'b000000000000000001100111;
		16'b1110001010010010 : data_out =  24'b000000000000000001100111;
		16'b1110001010010100 : data_out =  24'b000000000000000001100111;
		16'b1110001010010110 : data_out =  24'b000000000000000001100111;
		16'b1110001010011000 : data_out =  24'b000000000000000001100111;
		16'b1110001010011010 : data_out =  24'b000000000000000001100111;
		16'b1110001010011100 : data_out =  24'b000000000000000001100111;
		16'b1110001010011110 : data_out =  24'b000000000000000001101000;
		16'b1110001010100000 : data_out =  24'b000000000000000001101000;
		16'b1110001010100010 : data_out =  24'b000000000000000001101000;
		16'b1110001010100100 : data_out =  24'b000000000000000001101000;
		16'b1110001010100110 : data_out =  24'b000000000000000001101000;
		16'b1110001010101000 : data_out =  24'b000000000000000001101000;
		16'b1110001010101010 : data_out =  24'b000000000000000001101000;
		16'b1110001010101101 : data_out =  24'b000000000000000001101000;
		16'b1110001010101111 : data_out =  24'b000000000000000001101000;
		16'b1110001010110001 : data_out =  24'b000000000000000001101000;
		16'b1110001010110011 : data_out =  24'b000000000000000001101001;
		16'b1110001010110101 : data_out =  24'b000000000000000001101001;
		16'b1110001010110111 : data_out =  24'b000000000000000001101001;
		16'b1110001010111001 : data_out =  24'b000000000000000001101001;
		16'b1110001010111011 : data_out =  24'b000000000000000001101001;
		16'b1110001010111101 : data_out =  24'b000000000000000001101001;
		16'b1110001010111111 : data_out =  24'b000000000000000001101001;
		16'b1110001011000001 : data_out =  24'b000000000000000001101001;
		16'b1110001011000011 : data_out =  24'b000000000000000001101001;
		16'b1110001011000101 : data_out =  24'b000000000000000001101010;
		16'b1110001011000111 : data_out =  24'b000000000000000001101010;
		16'b1110001011001001 : data_out =  24'b000000000000000001101010;
		16'b1110001011001011 : data_out =  24'b000000000000000001101010;
		16'b1110001011001101 : data_out =  24'b000000000000000001101010;
		16'b1110001011001111 : data_out =  24'b000000000000000001101010;
		16'b1110001011010001 : data_out =  24'b000000000000000001101010;
		16'b1110001011010011 : data_out =  24'b000000000000000001101010;
		16'b1110001011010101 : data_out =  24'b000000000000000001101010;
		16'b1110001011011000 : data_out =  24'b000000000000000001101010;
		16'b1110001011011010 : data_out =  24'b000000000000000001101011;
		16'b1110001011011100 : data_out =  24'b000000000000000001101011;
		16'b1110001011011110 : data_out =  24'b000000000000000001101011;
		16'b1110001011100000 : data_out =  24'b000000000000000001101011;
		16'b1110001011100010 : data_out =  24'b000000000000000001101011;
		16'b1110001011100100 : data_out =  24'b000000000000000001101011;
		16'b1110001011100110 : data_out =  24'b000000000000000001101011;
		16'b1110001011101000 : data_out =  24'b000000000000000001101011;
		16'b1110001011101010 : data_out =  24'b000000000000000001101011;
		16'b1110001011101100 : data_out =  24'b000000000000000001101100;
		16'b1110001011101110 : data_out =  24'b000000000000000001101100;
		16'b1110001011110000 : data_out =  24'b000000000000000001101100;
		16'b1110001011110010 : data_out =  24'b000000000000000001101100;
		16'b1110001011110100 : data_out =  24'b000000000000000001101100;
		16'b1110001011110110 : data_out =  24'b000000000000000001101100;
		16'b1110001011111000 : data_out =  24'b000000000000000001101100;
		16'b1110001011111010 : data_out =  24'b000000000000000001101100;
		16'b1110001011111100 : data_out =  24'b000000000000000001101100;
		16'b1110001011111110 : data_out =  24'b000000000000000001101101;
		16'b1110001100000001 : data_out =  24'b000000000000000001101101;
		16'b1110001100000011 : data_out =  24'b000000000000000001101101;
		16'b1110001100000101 : data_out =  24'b000000000000000001101101;
		16'b1110001100000111 : data_out =  24'b000000000000000001101101;
		16'b1110001100001001 : data_out =  24'b000000000000000001101101;
		16'b1110001100001011 : data_out =  24'b000000000000000001101101;
		16'b1110001100001101 : data_out =  24'b000000000000000001101101;
		16'b1110001100001111 : data_out =  24'b000000000000000001101101;
		16'b1110001100010001 : data_out =  24'b000000000000000001101110;
		16'b1110001100010011 : data_out =  24'b000000000000000001101110;
		16'b1110001100010101 : data_out =  24'b000000000000000001101110;
		16'b1110001100010111 : data_out =  24'b000000000000000001101110;
		16'b1110001100011001 : data_out =  24'b000000000000000001101110;
		16'b1110001100011011 : data_out =  24'b000000000000000001101110;
		16'b1110001100011101 : data_out =  24'b000000000000000001101110;
		16'b1110001100011111 : data_out =  24'b000000000000000001101110;
		16'b1110001100100001 : data_out =  24'b000000000000000001101110;
		16'b1110001100100011 : data_out =  24'b000000000000000001101111;
		16'b1110001100100101 : data_out =  24'b000000000000000001101111;
		16'b1110001100100111 : data_out =  24'b000000000000000001101111;
		16'b1110001100101001 : data_out =  24'b000000000000000001101111;
		16'b1110001100101100 : data_out =  24'b000000000000000001101111;
		16'b1110001100101110 : data_out =  24'b000000000000000001101111;
		16'b1110001100110000 : data_out =  24'b000000000000000001101111;
		16'b1110001100110010 : data_out =  24'b000000000000000001101111;
		16'b1110001100110100 : data_out =  24'b000000000000000001101111;
		16'b1110001100110110 : data_out =  24'b000000000000000001110000;
		16'b1110001100111000 : data_out =  24'b000000000000000001110000;
		16'b1110001100111010 : data_out =  24'b000000000000000001110000;
		16'b1110001100111100 : data_out =  24'b000000000000000001110000;
		16'b1110001100111110 : data_out =  24'b000000000000000001110000;
		16'b1110001101000000 : data_out =  24'b000000000000000001110000;
		16'b1110001101000010 : data_out =  24'b000000000000000001110000;
		16'b1110001101000100 : data_out =  24'b000000000000000001110000;
		16'b1110001101000110 : data_out =  24'b000000000000000001110000;
		16'b1110001101001000 : data_out =  24'b000000000000000001110001;
		16'b1110001101001010 : data_out =  24'b000000000000000001110001;
		16'b1110001101001100 : data_out =  24'b000000000000000001110001;
		16'b1110001101001110 : data_out =  24'b000000000000000001110001;
		16'b1110001101010000 : data_out =  24'b000000000000000001110001;
		16'b1110001101010010 : data_out =  24'b000000000000000001110001;
		16'b1110001101010100 : data_out =  24'b000000000000000001110001;
		16'b1110001101010111 : data_out =  24'b000000000000000001110001;
		16'b1110001101011001 : data_out =  24'b000000000000000001110001;
		16'b1110001101011011 : data_out =  24'b000000000000000001110010;
		16'b1110001101011101 : data_out =  24'b000000000000000001110010;
		16'b1110001101011111 : data_out =  24'b000000000000000001110010;
		16'b1110001101100001 : data_out =  24'b000000000000000001110010;
		16'b1110001101100011 : data_out =  24'b000000000000000001110010;
		16'b1110001101100101 : data_out =  24'b000000000000000001110010;
		16'b1110001101100111 : data_out =  24'b000000000000000001110010;
		16'b1110001101101001 : data_out =  24'b000000000000000001110010;
		16'b1110001101101011 : data_out =  24'b000000000000000001110010;
		16'b1110001101101101 : data_out =  24'b000000000000000001110011;
		16'b1110001101101111 : data_out =  24'b000000000000000001110011;
		16'b1110001101110001 : data_out =  24'b000000000000000001110011;
		16'b1110001101110011 : data_out =  24'b000000000000000001110011;
		16'b1110001101110101 : data_out =  24'b000000000000000001110011;
		16'b1110001101110111 : data_out =  24'b000000000000000001110011;
		16'b1110001101111001 : data_out =  24'b000000000000000001110011;
		16'b1110001101111011 : data_out =  24'b000000000000000001110011;
		16'b1110001101111101 : data_out =  24'b000000000000000001110100;
		16'b1110001101111111 : data_out =  24'b000000000000000001110100;
		16'b1110001110000010 : data_out =  24'b000000000000000001110100;
		16'b1110001110000100 : data_out =  24'b000000000000000001110100;
		16'b1110001110000110 : data_out =  24'b000000000000000001110100;
		16'b1110001110001000 : data_out =  24'b000000000000000001110100;
		16'b1110001110001010 : data_out =  24'b000000000000000001110100;
		16'b1110001110001100 : data_out =  24'b000000000000000001110100;
		16'b1110001110001110 : data_out =  24'b000000000000000001110100;
		16'b1110001110010000 : data_out =  24'b000000000000000001110101;
		16'b1110001110010010 : data_out =  24'b000000000000000001110101;
		16'b1110001110010100 : data_out =  24'b000000000000000001110101;
		16'b1110001110010110 : data_out =  24'b000000000000000001110101;
		16'b1110001110011000 : data_out =  24'b000000000000000001110101;
		16'b1110001110011010 : data_out =  24'b000000000000000001110101;
		16'b1110001110011100 : data_out =  24'b000000000000000001110101;
		16'b1110001110011110 : data_out =  24'b000000000000000001110101;
		16'b1110001110100000 : data_out =  24'b000000000000000001110110;
		16'b1110001110100010 : data_out =  24'b000000000000000001110110;
		16'b1110001110100100 : data_out =  24'b000000000000000001110110;
		16'b1110001110100110 : data_out =  24'b000000000000000001110110;
		16'b1110001110101000 : data_out =  24'b000000000000000001110110;
		16'b1110001110101010 : data_out =  24'b000000000000000001110110;
		16'b1110001110101101 : data_out =  24'b000000000000000001110110;
		16'b1110001110101111 : data_out =  24'b000000000000000001110110;
		16'b1110001110110001 : data_out =  24'b000000000000000001110110;
		16'b1110001110110011 : data_out =  24'b000000000000000001110111;
		16'b1110001110110101 : data_out =  24'b000000000000000001110111;
		16'b1110001110110111 : data_out =  24'b000000000000000001110111;
		16'b1110001110111001 : data_out =  24'b000000000000000001110111;
		16'b1110001110111011 : data_out =  24'b000000000000000001110111;
		16'b1110001110111101 : data_out =  24'b000000000000000001110111;
		16'b1110001110111111 : data_out =  24'b000000000000000001110111;
		16'b1110001111000001 : data_out =  24'b000000000000000001110111;
		16'b1110001111000011 : data_out =  24'b000000000000000001111000;
		16'b1110001111000101 : data_out =  24'b000000000000000001111000;
		16'b1110001111000111 : data_out =  24'b000000000000000001111000;
		16'b1110001111001001 : data_out =  24'b000000000000000001111000;
		16'b1110001111001011 : data_out =  24'b000000000000000001111000;
		16'b1110001111001101 : data_out =  24'b000000000000000001111000;
		16'b1110001111001111 : data_out =  24'b000000000000000001111000;
		16'b1110001111010001 : data_out =  24'b000000000000000001111000;
		16'b1110001111010011 : data_out =  24'b000000000000000001111000;
		16'b1110001111010101 : data_out =  24'b000000000000000001111001;
		16'b1110001111011000 : data_out =  24'b000000000000000001111001;
		16'b1110001111011010 : data_out =  24'b000000000000000001111001;
		16'b1110001111011100 : data_out =  24'b000000000000000001111001;
		16'b1110001111011110 : data_out =  24'b000000000000000001111001;
		16'b1110001111100000 : data_out =  24'b000000000000000001111001;
		16'b1110001111100010 : data_out =  24'b000000000000000001111001;
		16'b1110001111100100 : data_out =  24'b000000000000000001111001;
		16'b1110001111100110 : data_out =  24'b000000000000000001111010;
		16'b1110001111101000 : data_out =  24'b000000000000000001111010;
		16'b1110001111101010 : data_out =  24'b000000000000000001111010;
		16'b1110001111101100 : data_out =  24'b000000000000000001111010;
		16'b1110001111101110 : data_out =  24'b000000000000000001111010;
		16'b1110001111110000 : data_out =  24'b000000000000000001111010;
		16'b1110001111110010 : data_out =  24'b000000000000000001111010;
		16'b1110001111110100 : data_out =  24'b000000000000000001111010;
		16'b1110001111110110 : data_out =  24'b000000000000000001111011;
		16'b1110001111111000 : data_out =  24'b000000000000000001111011;
		16'b1110001111111010 : data_out =  24'b000000000000000001111011;
		16'b1110001111111100 : data_out =  24'b000000000000000001111011;
		16'b1110001111111110 : data_out =  24'b000000000000000001111011;
		16'b1110010000000001 : data_out =  24'b000000000000000001111011;
		16'b1110010000000011 : data_out =  24'b000000000000000001111011;
		16'b1110010000000101 : data_out =  24'b000000000000000001111011;
		16'b1110010000000111 : data_out =  24'b000000000000000001111100;
		16'b1110010000001001 : data_out =  24'b000000000000000001111100;
		16'b1110010000001011 : data_out =  24'b000000000000000001111100;
		16'b1110010000001101 : data_out =  24'b000000000000000001111100;
		16'b1110010000001111 : data_out =  24'b000000000000000001111100;
		16'b1110010000010001 : data_out =  24'b000000000000000001111100;
		16'b1110010000010011 : data_out =  24'b000000000000000001111100;
		16'b1110010000010101 : data_out =  24'b000000000000000001111100;
		16'b1110010000010111 : data_out =  24'b000000000000000001111101;
		16'b1110010000011001 : data_out =  24'b000000000000000001111101;
		16'b1110010000011011 : data_out =  24'b000000000000000001111101;
		16'b1110010000011101 : data_out =  24'b000000000000000001111101;
		16'b1110010000011111 : data_out =  24'b000000000000000001111101;
		16'b1110010000100001 : data_out =  24'b000000000000000001111101;
		16'b1110010000100011 : data_out =  24'b000000000000000001111101;
		16'b1110010000100101 : data_out =  24'b000000000000000001111101;
		16'b1110010000100111 : data_out =  24'b000000000000000001111110;
		16'b1110010000101001 : data_out =  24'b000000000000000001111110;
		16'b1110010000101100 : data_out =  24'b000000000000000001111110;
		16'b1110010000101110 : data_out =  24'b000000000000000001111110;
		16'b1110010000110000 : data_out =  24'b000000000000000001111110;
		16'b1110010000110010 : data_out =  24'b000000000000000001111110;
		16'b1110010000110100 : data_out =  24'b000000000000000001111110;
		16'b1110010000110110 : data_out =  24'b000000000000000001111110;
		16'b1110010000111000 : data_out =  24'b000000000000000001111111;
		16'b1110010000111010 : data_out =  24'b000000000000000001111111;
		16'b1110010000111100 : data_out =  24'b000000000000000001111111;
		16'b1110010000111110 : data_out =  24'b000000000000000001111111;
		16'b1110010001000000 : data_out =  24'b000000000000000001111111;
		16'b1110010001000010 : data_out =  24'b000000000000000001111111;
		16'b1110010001000100 : data_out =  24'b000000000000000001111111;
		16'b1110010001000110 : data_out =  24'b000000000000000001111111;
		16'b1110010001001000 : data_out =  24'b000000000000000010000000;
		16'b1110010001001010 : data_out =  24'b000000000000000010000000;
		16'b1110010001001100 : data_out =  24'b000000000000000010000000;
		16'b1110010001001110 : data_out =  24'b000000000000000010000000;
		16'b1110010001010000 : data_out =  24'b000000000000000010000000;
		16'b1110010001010010 : data_out =  24'b000000000000000010000000;
		16'b1110010001010100 : data_out =  24'b000000000000000010000000;
		16'b1110010001010111 : data_out =  24'b000000000000000010000000;
		16'b1110010001011001 : data_out =  24'b000000000000000010000001;
		16'b1110010001011011 : data_out =  24'b000000000000000010000001;
		16'b1110010001011101 : data_out =  24'b000000000000000010000001;
		16'b1110010001011111 : data_out =  24'b000000000000000010000001;
		16'b1110010001100001 : data_out =  24'b000000000000000010000001;
		16'b1110010001100011 : data_out =  24'b000000000000000010000001;
		16'b1110010001100101 : data_out =  24'b000000000000000010000001;
		16'b1110010001100111 : data_out =  24'b000000000000000010000010;
		16'b1110010001101001 : data_out =  24'b000000000000000010000010;
		16'b1110010001101011 : data_out =  24'b000000000000000010000010;
		16'b1110010001101101 : data_out =  24'b000000000000000010000010;
		16'b1110010001101111 : data_out =  24'b000000000000000010000010;
		16'b1110010001110001 : data_out =  24'b000000000000000010000010;
		16'b1110010001110011 : data_out =  24'b000000000000000010000010;
		16'b1110010001110101 : data_out =  24'b000000000000000010000010;
		16'b1110010001110111 : data_out =  24'b000000000000000010000011;
		16'b1110010001111001 : data_out =  24'b000000000000000010000011;
		16'b1110010001111011 : data_out =  24'b000000000000000010000011;
		16'b1110010001111101 : data_out =  24'b000000000000000010000011;
		16'b1110010001111111 : data_out =  24'b000000000000000010000011;
		16'b1110010010000010 : data_out =  24'b000000000000000010000011;
		16'b1110010010000100 : data_out =  24'b000000000000000010000011;
		16'b1110010010000110 : data_out =  24'b000000000000000010000011;
		16'b1110010010001000 : data_out =  24'b000000000000000010000100;
		16'b1110010010001010 : data_out =  24'b000000000000000010000100;
		16'b1110010010001100 : data_out =  24'b000000000000000010000100;
		16'b1110010010001110 : data_out =  24'b000000000000000010000100;
		16'b1110010010010000 : data_out =  24'b000000000000000010000100;
		16'b1110010010010010 : data_out =  24'b000000000000000010000100;
		16'b1110010010010100 : data_out =  24'b000000000000000010000100;
		16'b1110010010010110 : data_out =  24'b000000000000000010000101;
		16'b1110010010011000 : data_out =  24'b000000000000000010000101;
		16'b1110010010011010 : data_out =  24'b000000000000000010000101;
		16'b1110010010011100 : data_out =  24'b000000000000000010000101;
		16'b1110010010011110 : data_out =  24'b000000000000000010000101;
		16'b1110010010100000 : data_out =  24'b000000000000000010000101;
		16'b1110010010100010 : data_out =  24'b000000000000000010000101;
		16'b1110010010100100 : data_out =  24'b000000000000000010000101;
		16'b1110010010100110 : data_out =  24'b000000000000000010000110;
		16'b1110010010101000 : data_out =  24'b000000000000000010000110;
		16'b1110010010101010 : data_out =  24'b000000000000000010000110;
		16'b1110010010101101 : data_out =  24'b000000000000000010000110;
		16'b1110010010101111 : data_out =  24'b000000000000000010000110;
		16'b1110010010110001 : data_out =  24'b000000000000000010000110;
		16'b1110010010110011 : data_out =  24'b000000000000000010000110;
		16'b1110010010110101 : data_out =  24'b000000000000000010000111;
		16'b1110010010110111 : data_out =  24'b000000000000000010000111;
		16'b1110010010111001 : data_out =  24'b000000000000000010000111;
		16'b1110010010111011 : data_out =  24'b000000000000000010000111;
		16'b1110010010111101 : data_out =  24'b000000000000000010000111;
		16'b1110010010111111 : data_out =  24'b000000000000000010000111;
		16'b1110010011000001 : data_out =  24'b000000000000000010000111;
		16'b1110010011000011 : data_out =  24'b000000000000000010001000;
		16'b1110010011000101 : data_out =  24'b000000000000000010001000;
		16'b1110010011000111 : data_out =  24'b000000000000000010001000;
		16'b1110010011001001 : data_out =  24'b000000000000000010001000;
		16'b1110010011001011 : data_out =  24'b000000000000000010001000;
		16'b1110010011001101 : data_out =  24'b000000000000000010001000;
		16'b1110010011001111 : data_out =  24'b000000000000000010001000;
		16'b1110010011010001 : data_out =  24'b000000000000000010001000;
		16'b1110010011010011 : data_out =  24'b000000000000000010001001;
		16'b1110010011010101 : data_out =  24'b000000000000000010001001;
		16'b1110010011011000 : data_out =  24'b000000000000000010001001;
		16'b1110010011011010 : data_out =  24'b000000000000000010001001;
		16'b1110010011011100 : data_out =  24'b000000000000000010001001;
		16'b1110010011011110 : data_out =  24'b000000000000000010001001;
		16'b1110010011100000 : data_out =  24'b000000000000000010001001;
		16'b1110010011100010 : data_out =  24'b000000000000000010001010;
		16'b1110010011100100 : data_out =  24'b000000000000000010001010;
		16'b1110010011100110 : data_out =  24'b000000000000000010001010;
		16'b1110010011101000 : data_out =  24'b000000000000000010001010;
		16'b1110010011101010 : data_out =  24'b000000000000000010001010;
		16'b1110010011101100 : data_out =  24'b000000000000000010001010;
		16'b1110010011101110 : data_out =  24'b000000000000000010001010;
		16'b1110010011110000 : data_out =  24'b000000000000000010001011;
		16'b1110010011110010 : data_out =  24'b000000000000000010001011;
		16'b1110010011110100 : data_out =  24'b000000000000000010001011;
		16'b1110010011110110 : data_out =  24'b000000000000000010001011;
		16'b1110010011111000 : data_out =  24'b000000000000000010001011;
		16'b1110010011111010 : data_out =  24'b000000000000000010001011;
		16'b1110010011111100 : data_out =  24'b000000000000000010001011;
		16'b1110010011111110 : data_out =  24'b000000000000000010001100;
		16'b1110010100000001 : data_out =  24'b000000000000000010001100;
		16'b1110010100000011 : data_out =  24'b000000000000000010001100;
		16'b1110010100000101 : data_out =  24'b000000000000000010001100;
		16'b1110010100000111 : data_out =  24'b000000000000000010001100;
		16'b1110010100001001 : data_out =  24'b000000000000000010001100;
		16'b1110010100001011 : data_out =  24'b000000000000000010001100;
		16'b1110010100001101 : data_out =  24'b000000000000000010001101;
		16'b1110010100001111 : data_out =  24'b000000000000000010001101;
		16'b1110010100010001 : data_out =  24'b000000000000000010001101;
		16'b1110010100010011 : data_out =  24'b000000000000000010001101;
		16'b1110010100010101 : data_out =  24'b000000000000000010001101;
		16'b1110010100010111 : data_out =  24'b000000000000000010001101;
		16'b1110010100011001 : data_out =  24'b000000000000000010001101;
		16'b1110010100011011 : data_out =  24'b000000000000000010001101;
		16'b1110010100011101 : data_out =  24'b000000000000000010001110;
		16'b1110010100011111 : data_out =  24'b000000000000000010001110;
		16'b1110010100100001 : data_out =  24'b000000000000000010001110;
		16'b1110010100100011 : data_out =  24'b000000000000000010001110;
		16'b1110010100100101 : data_out =  24'b000000000000000010001110;
		16'b1110010100100111 : data_out =  24'b000000000000000010001110;
		16'b1110010100101001 : data_out =  24'b000000000000000010001110;
		16'b1110010100101100 : data_out =  24'b000000000000000010001111;
		16'b1110010100101110 : data_out =  24'b000000000000000010001111;
		16'b1110010100110000 : data_out =  24'b000000000000000010001111;
		16'b1110010100110010 : data_out =  24'b000000000000000010001111;
		16'b1110010100110100 : data_out =  24'b000000000000000010001111;
		16'b1110010100110110 : data_out =  24'b000000000000000010001111;
		16'b1110010100111000 : data_out =  24'b000000000000000010001111;
		16'b1110010100111010 : data_out =  24'b000000000000000010010000;
		16'b1110010100111100 : data_out =  24'b000000000000000010010000;
		16'b1110010100111110 : data_out =  24'b000000000000000010010000;
		16'b1110010101000000 : data_out =  24'b000000000000000010010000;
		16'b1110010101000010 : data_out =  24'b000000000000000010010000;
		16'b1110010101000100 : data_out =  24'b000000000000000010010000;
		16'b1110010101000110 : data_out =  24'b000000000000000010010001;
		16'b1110010101001000 : data_out =  24'b000000000000000010010001;
		16'b1110010101001010 : data_out =  24'b000000000000000010010001;
		16'b1110010101001100 : data_out =  24'b000000000000000010010001;
		16'b1110010101001110 : data_out =  24'b000000000000000010010001;
		16'b1110010101010000 : data_out =  24'b000000000000000010010001;
		16'b1110010101010010 : data_out =  24'b000000000000000010010001;
		16'b1110010101010100 : data_out =  24'b000000000000000010010010;
		16'b1110010101010111 : data_out =  24'b000000000000000010010010;
		16'b1110010101011001 : data_out =  24'b000000000000000010010010;
		16'b1110010101011011 : data_out =  24'b000000000000000010010010;
		16'b1110010101011101 : data_out =  24'b000000000000000010010010;
		16'b1110010101011111 : data_out =  24'b000000000000000010010010;
		16'b1110010101100001 : data_out =  24'b000000000000000010010010;
		16'b1110010101100011 : data_out =  24'b000000000000000010010011;
		16'b1110010101100101 : data_out =  24'b000000000000000010010011;
		16'b1110010101100111 : data_out =  24'b000000000000000010010011;
		16'b1110010101101001 : data_out =  24'b000000000000000010010011;
		16'b1110010101101011 : data_out =  24'b000000000000000010010011;
		16'b1110010101101101 : data_out =  24'b000000000000000010010011;
		16'b1110010101101111 : data_out =  24'b000000000000000010010011;
		16'b1110010101110001 : data_out =  24'b000000000000000010010100;
		16'b1110010101110011 : data_out =  24'b000000000000000010010100;
		16'b1110010101110101 : data_out =  24'b000000000000000010010100;
		16'b1110010101110111 : data_out =  24'b000000000000000010010100;
		16'b1110010101111001 : data_out =  24'b000000000000000010010100;
		16'b1110010101111011 : data_out =  24'b000000000000000010010100;
		16'b1110010101111101 : data_out =  24'b000000000000000010010100;
		16'b1110010101111111 : data_out =  24'b000000000000000010010101;
		16'b1110010110000010 : data_out =  24'b000000000000000010010101;
		16'b1110010110000100 : data_out =  24'b000000000000000010010101;
		16'b1110010110000110 : data_out =  24'b000000000000000010010101;
		16'b1110010110001000 : data_out =  24'b000000000000000010010101;
		16'b1110010110001010 : data_out =  24'b000000000000000010010101;
		16'b1110010110001100 : data_out =  24'b000000000000000010010110;
		16'b1110010110001110 : data_out =  24'b000000000000000010010110;
		16'b1110010110010000 : data_out =  24'b000000000000000010010110;
		16'b1110010110010010 : data_out =  24'b000000000000000010010110;
		16'b1110010110010100 : data_out =  24'b000000000000000010010110;
		16'b1110010110010110 : data_out =  24'b000000000000000010010110;
		16'b1110010110011000 : data_out =  24'b000000000000000010010110;
		16'b1110010110011010 : data_out =  24'b000000000000000010010111;
		16'b1110010110011100 : data_out =  24'b000000000000000010010111;
		16'b1110010110011110 : data_out =  24'b000000000000000010010111;
		16'b1110010110100000 : data_out =  24'b000000000000000010010111;
		16'b1110010110100010 : data_out =  24'b000000000000000010010111;
		16'b1110010110100100 : data_out =  24'b000000000000000010010111;
		16'b1110010110100110 : data_out =  24'b000000000000000010010111;
		16'b1110010110101000 : data_out =  24'b000000000000000010011000;
		16'b1110010110101010 : data_out =  24'b000000000000000010011000;
		16'b1110010110101101 : data_out =  24'b000000000000000010011000;
		16'b1110010110101111 : data_out =  24'b000000000000000010011000;
		16'b1110010110110001 : data_out =  24'b000000000000000010011000;
		16'b1110010110110011 : data_out =  24'b000000000000000010011000;
		16'b1110010110110101 : data_out =  24'b000000000000000010011001;
		16'b1110010110110111 : data_out =  24'b000000000000000010011001;
		16'b1110010110111001 : data_out =  24'b000000000000000010011001;
		16'b1110010110111011 : data_out =  24'b000000000000000010011001;
		16'b1110010110111101 : data_out =  24'b000000000000000010011001;
		16'b1110010110111111 : data_out =  24'b000000000000000010011001;
		16'b1110010111000001 : data_out =  24'b000000000000000010011001;
		16'b1110010111000011 : data_out =  24'b000000000000000010011010;
		16'b1110010111000101 : data_out =  24'b000000000000000010011010;
		16'b1110010111000111 : data_out =  24'b000000000000000010011010;
		16'b1110010111001001 : data_out =  24'b000000000000000010011010;
		16'b1110010111001011 : data_out =  24'b000000000000000010011010;
		16'b1110010111001101 : data_out =  24'b000000000000000010011010;
		16'b1110010111001111 : data_out =  24'b000000000000000010011011;
		16'b1110010111010001 : data_out =  24'b000000000000000010011011;
		16'b1110010111010011 : data_out =  24'b000000000000000010011011;
		16'b1110010111010101 : data_out =  24'b000000000000000010011011;
		16'b1110010111011000 : data_out =  24'b000000000000000010011011;
		16'b1110010111011010 : data_out =  24'b000000000000000010011011;
		16'b1110010111011100 : data_out =  24'b000000000000000010011011;
		16'b1110010111011110 : data_out =  24'b000000000000000010011100;
		16'b1110010111100000 : data_out =  24'b000000000000000010011100;
		16'b1110010111100010 : data_out =  24'b000000000000000010011100;
		16'b1110010111100100 : data_out =  24'b000000000000000010011100;
		16'b1110010111100110 : data_out =  24'b000000000000000010011100;
		16'b1110010111101000 : data_out =  24'b000000000000000010011100;
		16'b1110010111101010 : data_out =  24'b000000000000000010011101;
		16'b1110010111101100 : data_out =  24'b000000000000000010011101;
		16'b1110010111101110 : data_out =  24'b000000000000000010011101;
		16'b1110010111110000 : data_out =  24'b000000000000000010011101;
		16'b1110010111110010 : data_out =  24'b000000000000000010011101;
		16'b1110010111110100 : data_out =  24'b000000000000000010011101;
		16'b1110010111110110 : data_out =  24'b000000000000000010011110;
		16'b1110010111111000 : data_out =  24'b000000000000000010011110;
		16'b1110010111111010 : data_out =  24'b000000000000000010011110;
		16'b1110010111111100 : data_out =  24'b000000000000000010011110;
		16'b1110010111111110 : data_out =  24'b000000000000000010011110;
		16'b1110011000000001 : data_out =  24'b000000000000000010011110;
		16'b1110011000000011 : data_out =  24'b000000000000000010011110;
		16'b1110011000000101 : data_out =  24'b000000000000000010011111;
		16'b1110011000000111 : data_out =  24'b000000000000000010011111;
		16'b1110011000001001 : data_out =  24'b000000000000000010011111;
		16'b1110011000001011 : data_out =  24'b000000000000000010011111;
		16'b1110011000001101 : data_out =  24'b000000000000000010011111;
		16'b1110011000001111 : data_out =  24'b000000000000000010011111;
		16'b1110011000010001 : data_out =  24'b000000000000000010100000;
		16'b1110011000010011 : data_out =  24'b000000000000000010100000;
		16'b1110011000010101 : data_out =  24'b000000000000000010100000;
		16'b1110011000010111 : data_out =  24'b000000000000000010100000;
		16'b1110011000011001 : data_out =  24'b000000000000000010100000;
		16'b1110011000011011 : data_out =  24'b000000000000000010100000;
		16'b1110011000011101 : data_out =  24'b000000000000000010100001;
		16'b1110011000011111 : data_out =  24'b000000000000000010100001;
		16'b1110011000100001 : data_out =  24'b000000000000000010100001;
		16'b1110011000100011 : data_out =  24'b000000000000000010100001;
		16'b1110011000100101 : data_out =  24'b000000000000000010100001;
		16'b1110011000100111 : data_out =  24'b000000000000000010100001;
		16'b1110011000101001 : data_out =  24'b000000000000000010100010;
		16'b1110011000101100 : data_out =  24'b000000000000000010100010;
		16'b1110011000101110 : data_out =  24'b000000000000000010100010;
		16'b1110011000110000 : data_out =  24'b000000000000000010100010;
		16'b1110011000110010 : data_out =  24'b000000000000000010100010;
		16'b1110011000110100 : data_out =  24'b000000000000000010100010;
		16'b1110011000110110 : data_out =  24'b000000000000000010100011;
		16'b1110011000111000 : data_out =  24'b000000000000000010100011;
		16'b1110011000111010 : data_out =  24'b000000000000000010100011;
		16'b1110011000111100 : data_out =  24'b000000000000000010100011;
		16'b1110011000111110 : data_out =  24'b000000000000000010100011;
		16'b1110011001000000 : data_out =  24'b000000000000000010100011;
		16'b1110011001000010 : data_out =  24'b000000000000000010100011;
		16'b1110011001000100 : data_out =  24'b000000000000000010100100;
		16'b1110011001000110 : data_out =  24'b000000000000000010100100;
		16'b1110011001001000 : data_out =  24'b000000000000000010100100;
		16'b1110011001001010 : data_out =  24'b000000000000000010100100;
		16'b1110011001001100 : data_out =  24'b000000000000000010100100;
		16'b1110011001001110 : data_out =  24'b000000000000000010100100;
		16'b1110011001010000 : data_out =  24'b000000000000000010100101;
		16'b1110011001010010 : data_out =  24'b000000000000000010100101;
		16'b1110011001010100 : data_out =  24'b000000000000000010100101;
		16'b1110011001010111 : data_out =  24'b000000000000000010100101;
		16'b1110011001011001 : data_out =  24'b000000000000000010100101;
		16'b1110011001011011 : data_out =  24'b000000000000000010100101;
		16'b1110011001011101 : data_out =  24'b000000000000000010100110;
		16'b1110011001011111 : data_out =  24'b000000000000000010100110;
		16'b1110011001100001 : data_out =  24'b000000000000000010100110;
		16'b1110011001100011 : data_out =  24'b000000000000000010100110;
		16'b1110011001100101 : data_out =  24'b000000000000000010100110;
		16'b1110011001100111 : data_out =  24'b000000000000000010100110;
		16'b1110011001101001 : data_out =  24'b000000000000000010100111;
		16'b1110011001101011 : data_out =  24'b000000000000000010100111;
		16'b1110011001101101 : data_out =  24'b000000000000000010100111;
		16'b1110011001101111 : data_out =  24'b000000000000000010100111;
		16'b1110011001110001 : data_out =  24'b000000000000000010100111;
		16'b1110011001110011 : data_out =  24'b000000000000000010100111;
		16'b1110011001110101 : data_out =  24'b000000000000000010101000;
		16'b1110011001110111 : data_out =  24'b000000000000000010101000;
		16'b1110011001111001 : data_out =  24'b000000000000000010101000;
		16'b1110011001111011 : data_out =  24'b000000000000000010101000;
		16'b1110011001111101 : data_out =  24'b000000000000000010101000;
		16'b1110011001111111 : data_out =  24'b000000000000000010101000;
		16'b1110011010000010 : data_out =  24'b000000000000000010101001;
		16'b1110011010000100 : data_out =  24'b000000000000000010101001;
		16'b1110011010000110 : data_out =  24'b000000000000000010101001;
		16'b1110011010001000 : data_out =  24'b000000000000000010101001;
		16'b1110011010001010 : data_out =  24'b000000000000000010101001;
		16'b1110011010001100 : data_out =  24'b000000000000000010101001;
		16'b1110011010001110 : data_out =  24'b000000000000000010101010;
		16'b1110011010010000 : data_out =  24'b000000000000000010101010;
		16'b1110011010010010 : data_out =  24'b000000000000000010101010;
		16'b1110011010010100 : data_out =  24'b000000000000000010101010;
		16'b1110011010010110 : data_out =  24'b000000000000000010101010;
		16'b1110011010011000 : data_out =  24'b000000000000000010101011;
		16'b1110011010011010 : data_out =  24'b000000000000000010101011;
		16'b1110011010011100 : data_out =  24'b000000000000000010101011;
		16'b1110011010011110 : data_out =  24'b000000000000000010101011;
		16'b1110011010100000 : data_out =  24'b000000000000000010101011;
		16'b1110011010100010 : data_out =  24'b000000000000000010101011;
		16'b1110011010100100 : data_out =  24'b000000000000000010101100;
		16'b1110011010100110 : data_out =  24'b000000000000000010101100;
		16'b1110011010101000 : data_out =  24'b000000000000000010101100;
		16'b1110011010101010 : data_out =  24'b000000000000000010101100;
		16'b1110011010101101 : data_out =  24'b000000000000000010101100;
		16'b1110011010101111 : data_out =  24'b000000000000000010101100;
		16'b1110011010110001 : data_out =  24'b000000000000000010101101;
		16'b1110011010110011 : data_out =  24'b000000000000000010101101;
		16'b1110011010110101 : data_out =  24'b000000000000000010101101;
		16'b1110011010110111 : data_out =  24'b000000000000000010101101;
		16'b1110011010111001 : data_out =  24'b000000000000000010101101;
		16'b1110011010111011 : data_out =  24'b000000000000000010101101;
		16'b1110011010111101 : data_out =  24'b000000000000000010101110;
		16'b1110011010111111 : data_out =  24'b000000000000000010101110;
		16'b1110011011000001 : data_out =  24'b000000000000000010101110;
		16'b1110011011000011 : data_out =  24'b000000000000000010101110;
		16'b1110011011000101 : data_out =  24'b000000000000000010101110;
		16'b1110011011000111 : data_out =  24'b000000000000000010101110;
		16'b1110011011001001 : data_out =  24'b000000000000000010101111;
		16'b1110011011001011 : data_out =  24'b000000000000000010101111;
		16'b1110011011001101 : data_out =  24'b000000000000000010101111;
		16'b1110011011001111 : data_out =  24'b000000000000000010101111;
		16'b1110011011010001 : data_out =  24'b000000000000000010101111;
		16'b1110011011010011 : data_out =  24'b000000000000000010110000;
		16'b1110011011010101 : data_out =  24'b000000000000000010110000;
		16'b1110011011011000 : data_out =  24'b000000000000000010110000;
		16'b1110011011011010 : data_out =  24'b000000000000000010110000;
		16'b1110011011011100 : data_out =  24'b000000000000000010110000;
		16'b1110011011011110 : data_out =  24'b000000000000000010110000;
		16'b1110011011100000 : data_out =  24'b000000000000000010110001;
		16'b1110011011100010 : data_out =  24'b000000000000000010110001;
		16'b1110011011100100 : data_out =  24'b000000000000000010110001;
		16'b1110011011100110 : data_out =  24'b000000000000000010110001;
		16'b1110011011101000 : data_out =  24'b000000000000000010110001;
		16'b1110011011101010 : data_out =  24'b000000000000000010110001;
		16'b1110011011101100 : data_out =  24'b000000000000000010110010;
		16'b1110011011101110 : data_out =  24'b000000000000000010110010;
		16'b1110011011110000 : data_out =  24'b000000000000000010110010;
		16'b1110011011110010 : data_out =  24'b000000000000000010110010;
		16'b1110011011110100 : data_out =  24'b000000000000000010110010;
		16'b1110011011110110 : data_out =  24'b000000000000000010110011;
		16'b1110011011111000 : data_out =  24'b000000000000000010110011;
		16'b1110011011111010 : data_out =  24'b000000000000000010110011;
		16'b1110011011111100 : data_out =  24'b000000000000000010110011;
		16'b1110011011111110 : data_out =  24'b000000000000000010110011;
		16'b1110011100000001 : data_out =  24'b000000000000000010110011;
		16'b1110011100000011 : data_out =  24'b000000000000000010110100;
		16'b1110011100000101 : data_out =  24'b000000000000000010110100;
		16'b1110011100000111 : data_out =  24'b000000000000000010110100;
		16'b1110011100001001 : data_out =  24'b000000000000000010110100;
		16'b1110011100001011 : data_out =  24'b000000000000000010110100;
		16'b1110011100001101 : data_out =  24'b000000000000000010110101;
		16'b1110011100001111 : data_out =  24'b000000000000000010110101;
		16'b1110011100010001 : data_out =  24'b000000000000000010110101;
		16'b1110011100010011 : data_out =  24'b000000000000000010110101;
		16'b1110011100010101 : data_out =  24'b000000000000000010110101;
		16'b1110011100010111 : data_out =  24'b000000000000000010110101;
		16'b1110011100011001 : data_out =  24'b000000000000000010110110;
		16'b1110011100011011 : data_out =  24'b000000000000000010110110;
		16'b1110011100011101 : data_out =  24'b000000000000000010110110;
		16'b1110011100011111 : data_out =  24'b000000000000000010110110;
		16'b1110011100100001 : data_out =  24'b000000000000000010110110;
		16'b1110011100100011 : data_out =  24'b000000000000000010110111;
		16'b1110011100100101 : data_out =  24'b000000000000000010110111;
		16'b1110011100100111 : data_out =  24'b000000000000000010110111;
		16'b1110011100101001 : data_out =  24'b000000000000000010110111;
		16'b1110011100101100 : data_out =  24'b000000000000000010110111;
		16'b1110011100101110 : data_out =  24'b000000000000000010110111;
		16'b1110011100110000 : data_out =  24'b000000000000000010111000;
		16'b1110011100110010 : data_out =  24'b000000000000000010111000;
		16'b1110011100110100 : data_out =  24'b000000000000000010111000;
		16'b1110011100110110 : data_out =  24'b000000000000000010111000;
		16'b1110011100111000 : data_out =  24'b000000000000000010111000;
		16'b1110011100111010 : data_out =  24'b000000000000000010111001;
		16'b1110011100111100 : data_out =  24'b000000000000000010111001;
		16'b1110011100111110 : data_out =  24'b000000000000000010111001;
		16'b1110011101000000 : data_out =  24'b000000000000000010111001;
		16'b1110011101000010 : data_out =  24'b000000000000000010111001;
		16'b1110011101000100 : data_out =  24'b000000000000000010111010;
		16'b1110011101000110 : data_out =  24'b000000000000000010111010;
		16'b1110011101001000 : data_out =  24'b000000000000000010111010;
		16'b1110011101001010 : data_out =  24'b000000000000000010111010;
		16'b1110011101001100 : data_out =  24'b000000000000000010111010;
		16'b1110011101001110 : data_out =  24'b000000000000000010111010;
		16'b1110011101010000 : data_out =  24'b000000000000000010111011;
		16'b1110011101010010 : data_out =  24'b000000000000000010111011;
		16'b1110011101010100 : data_out =  24'b000000000000000010111011;
		16'b1110011101010111 : data_out =  24'b000000000000000010111011;
		16'b1110011101011001 : data_out =  24'b000000000000000010111011;
		16'b1110011101011011 : data_out =  24'b000000000000000010111100;
		16'b1110011101011101 : data_out =  24'b000000000000000010111100;
		16'b1110011101011111 : data_out =  24'b000000000000000010111100;
		16'b1110011101100001 : data_out =  24'b000000000000000010111100;
		16'b1110011101100011 : data_out =  24'b000000000000000010111100;
		16'b1110011101100101 : data_out =  24'b000000000000000010111101;
		16'b1110011101100111 : data_out =  24'b000000000000000010111101;
		16'b1110011101101001 : data_out =  24'b000000000000000010111101;
		16'b1110011101101011 : data_out =  24'b000000000000000010111101;
		16'b1110011101101101 : data_out =  24'b000000000000000010111101;
		16'b1110011101101111 : data_out =  24'b000000000000000010111101;
		16'b1110011101110001 : data_out =  24'b000000000000000010111110;
		16'b1110011101110011 : data_out =  24'b000000000000000010111110;
		16'b1110011101110101 : data_out =  24'b000000000000000010111110;
		16'b1110011101110111 : data_out =  24'b000000000000000010111110;
		16'b1110011101111001 : data_out =  24'b000000000000000010111110;
		16'b1110011101111011 : data_out =  24'b000000000000000010111111;
		16'b1110011101111101 : data_out =  24'b000000000000000010111111;
		16'b1110011101111111 : data_out =  24'b000000000000000010111111;
		16'b1110011110000010 : data_out =  24'b000000000000000010111111;
		16'b1110011110000100 : data_out =  24'b000000000000000010111111;
		16'b1110011110000110 : data_out =  24'b000000000000000011000000;
		16'b1110011110001000 : data_out =  24'b000000000000000011000000;
		16'b1110011110001010 : data_out =  24'b000000000000000011000000;
		16'b1110011110001100 : data_out =  24'b000000000000000011000000;
		16'b1110011110001110 : data_out =  24'b000000000000000011000000;
		16'b1110011110010000 : data_out =  24'b000000000000000011000001;
		16'b1110011110010010 : data_out =  24'b000000000000000011000001;
		16'b1110011110010100 : data_out =  24'b000000000000000011000001;
		16'b1110011110010110 : data_out =  24'b000000000000000011000001;
		16'b1110011110011000 : data_out =  24'b000000000000000011000001;
		16'b1110011110011010 : data_out =  24'b000000000000000011000001;
		16'b1110011110011100 : data_out =  24'b000000000000000011000010;
		16'b1110011110011110 : data_out =  24'b000000000000000011000010;
		16'b1110011110100000 : data_out =  24'b000000000000000011000010;
		16'b1110011110100010 : data_out =  24'b000000000000000011000010;
		16'b1110011110100100 : data_out =  24'b000000000000000011000010;
		16'b1110011110100110 : data_out =  24'b000000000000000011000011;
		16'b1110011110101000 : data_out =  24'b000000000000000011000011;
		16'b1110011110101010 : data_out =  24'b000000000000000011000011;
		16'b1110011110101101 : data_out =  24'b000000000000000011000011;
		16'b1110011110101111 : data_out =  24'b000000000000000011000011;
		16'b1110011110110001 : data_out =  24'b000000000000000011000100;
		16'b1110011110110011 : data_out =  24'b000000000000000011000100;
		16'b1110011110110101 : data_out =  24'b000000000000000011000100;
		16'b1110011110110111 : data_out =  24'b000000000000000011000100;
		16'b1110011110111001 : data_out =  24'b000000000000000011000100;
		16'b1110011110111011 : data_out =  24'b000000000000000011000101;
		16'b1110011110111101 : data_out =  24'b000000000000000011000101;
		16'b1110011110111111 : data_out =  24'b000000000000000011000101;
		16'b1110011111000001 : data_out =  24'b000000000000000011000101;
		16'b1110011111000011 : data_out =  24'b000000000000000011000101;
		16'b1110011111000101 : data_out =  24'b000000000000000011000110;
		16'b1110011111000111 : data_out =  24'b000000000000000011000110;
		16'b1110011111001001 : data_out =  24'b000000000000000011000110;
		16'b1110011111001011 : data_out =  24'b000000000000000011000110;
		16'b1110011111001101 : data_out =  24'b000000000000000011000110;
		16'b1110011111001111 : data_out =  24'b000000000000000011000111;
		16'b1110011111010001 : data_out =  24'b000000000000000011000111;
		16'b1110011111010011 : data_out =  24'b000000000000000011000111;
		16'b1110011111010101 : data_out =  24'b000000000000000011000111;
		16'b1110011111011000 : data_out =  24'b000000000000000011000111;
		16'b1110011111011010 : data_out =  24'b000000000000000011001000;
		16'b1110011111011100 : data_out =  24'b000000000000000011001000;
		16'b1110011111011110 : data_out =  24'b000000000000000011001000;
		16'b1110011111100000 : data_out =  24'b000000000000000011001000;
		16'b1110011111100010 : data_out =  24'b000000000000000011001000;
		16'b1110011111100100 : data_out =  24'b000000000000000011001001;
		16'b1110011111100110 : data_out =  24'b000000000000000011001001;
		16'b1110011111101000 : data_out =  24'b000000000000000011001001;
		16'b1110011111101010 : data_out =  24'b000000000000000011001001;
		16'b1110011111101100 : data_out =  24'b000000000000000011001001;
		16'b1110011111101110 : data_out =  24'b000000000000000011001010;
		16'b1110011111110000 : data_out =  24'b000000000000000011001010;
		16'b1110011111110010 : data_out =  24'b000000000000000011001010;
		16'b1110011111110100 : data_out =  24'b000000000000000011001010;
		16'b1110011111110110 : data_out =  24'b000000000000000011001010;
		16'b1110011111111000 : data_out =  24'b000000000000000011001011;
		16'b1110011111111010 : data_out =  24'b000000000000000011001011;
		16'b1110011111111100 : data_out =  24'b000000000000000011001011;
		16'b1110011111111110 : data_out =  24'b000000000000000011001011;
		16'b1110100000000001 : data_out =  24'b000000000000000011001011;
		16'b1110100000000011 : data_out =  24'b000000000000000011001100;
		16'b1110100000000101 : data_out =  24'b000000000000000011001100;
		16'b1110100000000111 : data_out =  24'b000000000000000011001100;
		16'b1110100000001001 : data_out =  24'b000000000000000011001100;
		16'b1110100000001011 : data_out =  24'b000000000000000011001100;
		16'b1110100000001101 : data_out =  24'b000000000000000011001101;
		16'b1110100000001111 : data_out =  24'b000000000000000011001101;
		16'b1110100000010001 : data_out =  24'b000000000000000011001101;
		16'b1110100000010011 : data_out =  24'b000000000000000011001101;
		16'b1110100000010101 : data_out =  24'b000000000000000011001101;
		16'b1110100000010111 : data_out =  24'b000000000000000011001110;
		16'b1110100000011001 : data_out =  24'b000000000000000011001110;
		16'b1110100000011011 : data_out =  24'b000000000000000011001110;
		16'b1110100000011101 : data_out =  24'b000000000000000011001110;
		16'b1110100000011111 : data_out =  24'b000000000000000011001111;
		16'b1110100000100001 : data_out =  24'b000000000000000011001111;
		16'b1110100000100011 : data_out =  24'b000000000000000011001111;
		16'b1110100000100101 : data_out =  24'b000000000000000011001111;
		16'b1110100000100111 : data_out =  24'b000000000000000011001111;
		16'b1110100000101001 : data_out =  24'b000000000000000011010000;
		16'b1110100000101100 : data_out =  24'b000000000000000011010000;
		16'b1110100000101110 : data_out =  24'b000000000000000011010000;
		16'b1110100000110000 : data_out =  24'b000000000000000011010000;
		16'b1110100000110010 : data_out =  24'b000000000000000011010000;
		16'b1110100000110100 : data_out =  24'b000000000000000011010001;
		16'b1110100000110110 : data_out =  24'b000000000000000011010001;
		16'b1110100000111000 : data_out =  24'b000000000000000011010001;
		16'b1110100000111010 : data_out =  24'b000000000000000011010001;
		16'b1110100000111100 : data_out =  24'b000000000000000011010001;
		16'b1110100000111110 : data_out =  24'b000000000000000011010010;
		16'b1110100001000000 : data_out =  24'b000000000000000011010010;
		16'b1110100001000010 : data_out =  24'b000000000000000011010010;
		16'b1110100001000100 : data_out =  24'b000000000000000011010010;
		16'b1110100001000110 : data_out =  24'b000000000000000011010010;
		16'b1110100001001000 : data_out =  24'b000000000000000011010011;
		16'b1110100001001010 : data_out =  24'b000000000000000011010011;
		16'b1110100001001100 : data_out =  24'b000000000000000011010011;
		16'b1110100001001110 : data_out =  24'b000000000000000011010011;
		16'b1110100001010000 : data_out =  24'b000000000000000011010100;
		16'b1110100001010010 : data_out =  24'b000000000000000011010100;
		16'b1110100001010100 : data_out =  24'b000000000000000011010100;
		16'b1110100001010111 : data_out =  24'b000000000000000011010100;
		16'b1110100001011001 : data_out =  24'b000000000000000011010100;
		16'b1110100001011011 : data_out =  24'b000000000000000011010101;
		16'b1110100001011101 : data_out =  24'b000000000000000011010101;
		16'b1110100001011111 : data_out =  24'b000000000000000011010101;
		16'b1110100001100001 : data_out =  24'b000000000000000011010101;
		16'b1110100001100011 : data_out =  24'b000000000000000011010101;
		16'b1110100001100101 : data_out =  24'b000000000000000011010110;
		16'b1110100001100111 : data_out =  24'b000000000000000011010110;
		16'b1110100001101001 : data_out =  24'b000000000000000011010110;
		16'b1110100001101011 : data_out =  24'b000000000000000011010110;
		16'b1110100001101101 : data_out =  24'b000000000000000011010111;
		16'b1110100001101111 : data_out =  24'b000000000000000011010111;
		16'b1110100001110001 : data_out =  24'b000000000000000011010111;
		16'b1110100001110011 : data_out =  24'b000000000000000011010111;
		16'b1110100001110101 : data_out =  24'b000000000000000011010111;
		16'b1110100001110111 : data_out =  24'b000000000000000011011000;
		16'b1110100001111001 : data_out =  24'b000000000000000011011000;
		16'b1110100001111011 : data_out =  24'b000000000000000011011000;
		16'b1110100001111101 : data_out =  24'b000000000000000011011000;
		16'b1110100001111111 : data_out =  24'b000000000000000011011000;
		16'b1110100010000010 : data_out =  24'b000000000000000011011001;
		16'b1110100010000100 : data_out =  24'b000000000000000011011001;
		16'b1110100010000110 : data_out =  24'b000000000000000011011001;
		16'b1110100010001000 : data_out =  24'b000000000000000011011001;
		16'b1110100010001010 : data_out =  24'b000000000000000011011010;
		16'b1110100010001100 : data_out =  24'b000000000000000011011010;
		16'b1110100010001110 : data_out =  24'b000000000000000011011010;
		16'b1110100010010000 : data_out =  24'b000000000000000011011010;
		16'b1110100010010010 : data_out =  24'b000000000000000011011010;
		16'b1110100010010100 : data_out =  24'b000000000000000011011011;
		16'b1110100010010110 : data_out =  24'b000000000000000011011011;
		16'b1110100010011000 : data_out =  24'b000000000000000011011011;
		16'b1110100010011010 : data_out =  24'b000000000000000011011011;
		16'b1110100010011100 : data_out =  24'b000000000000000011011100;
		16'b1110100010011110 : data_out =  24'b000000000000000011011100;
		16'b1110100010100000 : data_out =  24'b000000000000000011011100;
		16'b1110100010100010 : data_out =  24'b000000000000000011011100;
		16'b1110100010100100 : data_out =  24'b000000000000000011011100;
		16'b1110100010100110 : data_out =  24'b000000000000000011011101;
		16'b1110100010101000 : data_out =  24'b000000000000000011011101;
		16'b1110100010101010 : data_out =  24'b000000000000000011011101;
		16'b1110100010101101 : data_out =  24'b000000000000000011011101;
		16'b1110100010101111 : data_out =  24'b000000000000000011011110;
		16'b1110100010110001 : data_out =  24'b000000000000000011011110;
		16'b1110100010110011 : data_out =  24'b000000000000000011011110;
		16'b1110100010110101 : data_out =  24'b000000000000000011011110;
		16'b1110100010110111 : data_out =  24'b000000000000000011011110;
		16'b1110100010111001 : data_out =  24'b000000000000000011011111;
		16'b1110100010111011 : data_out =  24'b000000000000000011011111;
		16'b1110100010111101 : data_out =  24'b000000000000000011011111;
		16'b1110100010111111 : data_out =  24'b000000000000000011011111;
		16'b1110100011000001 : data_out =  24'b000000000000000011100000;
		16'b1110100011000011 : data_out =  24'b000000000000000011100000;
		16'b1110100011000101 : data_out =  24'b000000000000000011100000;
		16'b1110100011000111 : data_out =  24'b000000000000000011100000;
		16'b1110100011001001 : data_out =  24'b000000000000000011100000;
		16'b1110100011001011 : data_out =  24'b000000000000000011100001;
		16'b1110100011001101 : data_out =  24'b000000000000000011100001;
		16'b1110100011001111 : data_out =  24'b000000000000000011100001;
		16'b1110100011010001 : data_out =  24'b000000000000000011100001;
		16'b1110100011010011 : data_out =  24'b000000000000000011100010;
		16'b1110100011010101 : data_out =  24'b000000000000000011100010;
		16'b1110100011011000 : data_out =  24'b000000000000000011100010;
		16'b1110100011011010 : data_out =  24'b000000000000000011100010;
		16'b1110100011011100 : data_out =  24'b000000000000000011100010;
		16'b1110100011011110 : data_out =  24'b000000000000000011100011;
		16'b1110100011100000 : data_out =  24'b000000000000000011100011;
		16'b1110100011100010 : data_out =  24'b000000000000000011100011;
		16'b1110100011100100 : data_out =  24'b000000000000000011100011;
		16'b1110100011100110 : data_out =  24'b000000000000000011100100;
		16'b1110100011101000 : data_out =  24'b000000000000000011100100;
		16'b1110100011101010 : data_out =  24'b000000000000000011100100;
		16'b1110100011101100 : data_out =  24'b000000000000000011100100;
		16'b1110100011101110 : data_out =  24'b000000000000000011100101;
		16'b1110100011110000 : data_out =  24'b000000000000000011100101;
		16'b1110100011110010 : data_out =  24'b000000000000000011100101;
		16'b1110100011110100 : data_out =  24'b000000000000000011100101;
		16'b1110100011110110 : data_out =  24'b000000000000000011100101;
		16'b1110100011111000 : data_out =  24'b000000000000000011100110;
		16'b1110100011111010 : data_out =  24'b000000000000000011100110;
		16'b1110100011111100 : data_out =  24'b000000000000000011100110;
		16'b1110100011111110 : data_out =  24'b000000000000000011100110;
		16'b1110100100000001 : data_out =  24'b000000000000000011100111;
		16'b1110100100000011 : data_out =  24'b000000000000000011100111;
		16'b1110100100000101 : data_out =  24'b000000000000000011100111;
		16'b1110100100000111 : data_out =  24'b000000000000000011100111;
		16'b1110100100001001 : data_out =  24'b000000000000000011101000;
		16'b1110100100001011 : data_out =  24'b000000000000000011101000;
		16'b1110100100001101 : data_out =  24'b000000000000000011101000;
		16'b1110100100001111 : data_out =  24'b000000000000000011101000;
		16'b1110100100010001 : data_out =  24'b000000000000000011101000;
		16'b1110100100010011 : data_out =  24'b000000000000000011101001;
		16'b1110100100010101 : data_out =  24'b000000000000000011101001;
		16'b1110100100010111 : data_out =  24'b000000000000000011101001;
		16'b1110100100011001 : data_out =  24'b000000000000000011101001;
		16'b1110100100011011 : data_out =  24'b000000000000000011101010;
		16'b1110100100011101 : data_out =  24'b000000000000000011101010;
		16'b1110100100011111 : data_out =  24'b000000000000000011101010;
		16'b1110100100100001 : data_out =  24'b000000000000000011101010;
		16'b1110100100100011 : data_out =  24'b000000000000000011101011;
		16'b1110100100100101 : data_out =  24'b000000000000000011101011;
		16'b1110100100100111 : data_out =  24'b000000000000000011101011;
		16'b1110100100101001 : data_out =  24'b000000000000000011101011;
		16'b1110100100101100 : data_out =  24'b000000000000000011101011;
		16'b1110100100101110 : data_out =  24'b000000000000000011101100;
		16'b1110100100110000 : data_out =  24'b000000000000000011101100;
		16'b1110100100110010 : data_out =  24'b000000000000000011101100;
		16'b1110100100110100 : data_out =  24'b000000000000000011101100;
		16'b1110100100110110 : data_out =  24'b000000000000000011101101;
		16'b1110100100111000 : data_out =  24'b000000000000000011101101;
		16'b1110100100111010 : data_out =  24'b000000000000000011101101;
		16'b1110100100111100 : data_out =  24'b000000000000000011101101;
		16'b1110100100111110 : data_out =  24'b000000000000000011101110;
		16'b1110100101000000 : data_out =  24'b000000000000000011101110;
		16'b1110100101000010 : data_out =  24'b000000000000000011101110;
		16'b1110100101000100 : data_out =  24'b000000000000000011101110;
		16'b1110100101000110 : data_out =  24'b000000000000000011101111;
		16'b1110100101001000 : data_out =  24'b000000000000000011101111;
		16'b1110100101001010 : data_out =  24'b000000000000000011101111;
		16'b1110100101001100 : data_out =  24'b000000000000000011101111;
		16'b1110100101001110 : data_out =  24'b000000000000000011110000;
		16'b1110100101010000 : data_out =  24'b000000000000000011110000;
		16'b1110100101010010 : data_out =  24'b000000000000000011110000;
		16'b1110100101010100 : data_out =  24'b000000000000000011110000;
		16'b1110100101010111 : data_out =  24'b000000000000000011110000;
		16'b1110100101011001 : data_out =  24'b000000000000000011110001;
		16'b1110100101011011 : data_out =  24'b000000000000000011110001;
		16'b1110100101011101 : data_out =  24'b000000000000000011110001;
		16'b1110100101011111 : data_out =  24'b000000000000000011110001;
		16'b1110100101100001 : data_out =  24'b000000000000000011110010;
		16'b1110100101100011 : data_out =  24'b000000000000000011110010;
		16'b1110100101100101 : data_out =  24'b000000000000000011110010;
		16'b1110100101100111 : data_out =  24'b000000000000000011110010;
		16'b1110100101101001 : data_out =  24'b000000000000000011110011;
		16'b1110100101101011 : data_out =  24'b000000000000000011110011;
		16'b1110100101101101 : data_out =  24'b000000000000000011110011;
		16'b1110100101101111 : data_out =  24'b000000000000000011110011;
		16'b1110100101110001 : data_out =  24'b000000000000000011110100;
		16'b1110100101110011 : data_out =  24'b000000000000000011110100;
		16'b1110100101110101 : data_out =  24'b000000000000000011110100;
		16'b1110100101110111 : data_out =  24'b000000000000000011110100;
		16'b1110100101111001 : data_out =  24'b000000000000000011110101;
		16'b1110100101111011 : data_out =  24'b000000000000000011110101;
		16'b1110100101111101 : data_out =  24'b000000000000000011110101;
		16'b1110100101111111 : data_out =  24'b000000000000000011110101;
		16'b1110100110000010 : data_out =  24'b000000000000000011110110;
		16'b1110100110000100 : data_out =  24'b000000000000000011110110;
		16'b1110100110000110 : data_out =  24'b000000000000000011110110;
		16'b1110100110001000 : data_out =  24'b000000000000000011110110;
		16'b1110100110001010 : data_out =  24'b000000000000000011110111;
		16'b1110100110001100 : data_out =  24'b000000000000000011110111;
		16'b1110100110001110 : data_out =  24'b000000000000000011110111;
		16'b1110100110010000 : data_out =  24'b000000000000000011110111;
		16'b1110100110010010 : data_out =  24'b000000000000000011111000;
		16'b1110100110010100 : data_out =  24'b000000000000000011111000;
		16'b1110100110010110 : data_out =  24'b000000000000000011111000;
		16'b1110100110011000 : data_out =  24'b000000000000000011111000;
		16'b1110100110011010 : data_out =  24'b000000000000000011111001;
		16'b1110100110011100 : data_out =  24'b000000000000000011111001;
		16'b1110100110011110 : data_out =  24'b000000000000000011111001;
		16'b1110100110100000 : data_out =  24'b000000000000000011111001;
		16'b1110100110100010 : data_out =  24'b000000000000000011111010;
		16'b1110100110100100 : data_out =  24'b000000000000000011111010;
		16'b1110100110100110 : data_out =  24'b000000000000000011111010;
		16'b1110100110101000 : data_out =  24'b000000000000000011111010;
		16'b1110100110101010 : data_out =  24'b000000000000000011111011;
		16'b1110100110101101 : data_out =  24'b000000000000000011111011;
		16'b1110100110101111 : data_out =  24'b000000000000000011111011;
		16'b1110100110110001 : data_out =  24'b000000000000000011111011;
		16'b1110100110110011 : data_out =  24'b000000000000000011111100;
		16'b1110100110110101 : data_out =  24'b000000000000000011111100;
		16'b1110100110110111 : data_out =  24'b000000000000000011111100;
		16'b1110100110111001 : data_out =  24'b000000000000000011111100;
		16'b1110100110111011 : data_out =  24'b000000000000000011111101;
		16'b1110100110111101 : data_out =  24'b000000000000000011111101;
		16'b1110100110111111 : data_out =  24'b000000000000000011111101;
		16'b1110100111000001 : data_out =  24'b000000000000000011111101;
		16'b1110100111000011 : data_out =  24'b000000000000000011111110;
		16'b1110100111000101 : data_out =  24'b000000000000000011111110;
		16'b1110100111000111 : data_out =  24'b000000000000000011111110;
		16'b1110100111001001 : data_out =  24'b000000000000000011111110;
		16'b1110100111001011 : data_out =  24'b000000000000000011111111;
		16'b1110100111001101 : data_out =  24'b000000000000000011111111;
		16'b1110100111001111 : data_out =  24'b000000000000000011111111;
		16'b1110100111010001 : data_out =  24'b000000000000000011111111;
		16'b1110100111010011 : data_out =  24'b000000000000000100000000;
		16'b1110100111010101 : data_out =  24'b000000000000000100000000;
		16'b1110100111011000 : data_out =  24'b000000000000000100000000;
		16'b1110100111011010 : data_out =  24'b000000000000000100000000;
		16'b1110100111011100 : data_out =  24'b000000000000000100000001;
		16'b1110100111011110 : data_out =  24'b000000000000000100000001;
		16'b1110100111100000 : data_out =  24'b000000000000000100000001;
		16'b1110100111100010 : data_out =  24'b000000000000000100000001;
		16'b1110100111100100 : data_out =  24'b000000000000000100000010;
		16'b1110100111100110 : data_out =  24'b000000000000000100000010;
		16'b1110100111101000 : data_out =  24'b000000000000000100000010;
		16'b1110100111101010 : data_out =  24'b000000000000000100000010;
		16'b1110100111101100 : data_out =  24'b000000000000000100000011;
		16'b1110100111101110 : data_out =  24'b000000000000000100000011;
		16'b1110100111110000 : data_out =  24'b000000000000000100000011;
		16'b1110100111110010 : data_out =  24'b000000000000000100000100;
		16'b1110100111110100 : data_out =  24'b000000000000000100000100;
		16'b1110100111110110 : data_out =  24'b000000000000000100000100;
		16'b1110100111111000 : data_out =  24'b000000000000000100000100;
		16'b1110100111111010 : data_out =  24'b000000000000000100000101;
		16'b1110100111111100 : data_out =  24'b000000000000000100000101;
		16'b1110100111111110 : data_out =  24'b000000000000000100000101;
		16'b1110101000000001 : data_out =  24'b000000000000000100000101;
		16'b1110101000000011 : data_out =  24'b000000000000000100000110;
		16'b1110101000000101 : data_out =  24'b000000000000000100000110;
		16'b1110101000000111 : data_out =  24'b000000000000000100000110;
		16'b1110101000001001 : data_out =  24'b000000000000000100000110;
		16'b1110101000001011 : data_out =  24'b000000000000000100000111;
		16'b1110101000001101 : data_out =  24'b000000000000000100000111;
		16'b1110101000001111 : data_out =  24'b000000000000000100000111;
		16'b1110101000010001 : data_out =  24'b000000000000000100000111;
		16'b1110101000010011 : data_out =  24'b000000000000000100001000;
		16'b1110101000010101 : data_out =  24'b000000000000000100001000;
		16'b1110101000010111 : data_out =  24'b000000000000000100001000;
		16'b1110101000011001 : data_out =  24'b000000000000000100001001;
		16'b1110101000011011 : data_out =  24'b000000000000000100001001;
		16'b1110101000011101 : data_out =  24'b000000000000000100001001;
		16'b1110101000011111 : data_out =  24'b000000000000000100001001;
		16'b1110101000100001 : data_out =  24'b000000000000000100001010;
		16'b1110101000100011 : data_out =  24'b000000000000000100001010;
		16'b1110101000100101 : data_out =  24'b000000000000000100001010;
		16'b1110101000100111 : data_out =  24'b000000000000000100001010;
		16'b1110101000101001 : data_out =  24'b000000000000000100001011;
		16'b1110101000101100 : data_out =  24'b000000000000000100001011;
		16'b1110101000101110 : data_out =  24'b000000000000000100001011;
		16'b1110101000110000 : data_out =  24'b000000000000000100001011;
		16'b1110101000110010 : data_out =  24'b000000000000000100001100;
		16'b1110101000110100 : data_out =  24'b000000000000000100001100;
		16'b1110101000110110 : data_out =  24'b000000000000000100001100;
		16'b1110101000111000 : data_out =  24'b000000000000000100001101;
		16'b1110101000111010 : data_out =  24'b000000000000000100001101;
		16'b1110101000111100 : data_out =  24'b000000000000000100001101;
		16'b1110101000111110 : data_out =  24'b000000000000000100001101;
		16'b1110101001000000 : data_out =  24'b000000000000000100001110;
		16'b1110101001000010 : data_out =  24'b000000000000000100001110;
		16'b1110101001000100 : data_out =  24'b000000000000000100001110;
		16'b1110101001000110 : data_out =  24'b000000000000000100001110;
		16'b1110101001001000 : data_out =  24'b000000000000000100001111;
		16'b1110101001001010 : data_out =  24'b000000000000000100001111;
		16'b1110101001001100 : data_out =  24'b000000000000000100001111;
		16'b1110101001001110 : data_out =  24'b000000000000000100001111;
		16'b1110101001010000 : data_out =  24'b000000000000000100010000;
		16'b1110101001010010 : data_out =  24'b000000000000000100010000;
		16'b1110101001010100 : data_out =  24'b000000000000000100010000;
		16'b1110101001010111 : data_out =  24'b000000000000000100010001;
		16'b1110101001011001 : data_out =  24'b000000000000000100010001;
		16'b1110101001011011 : data_out =  24'b000000000000000100010001;
		16'b1110101001011101 : data_out =  24'b000000000000000100010001;
		16'b1110101001011111 : data_out =  24'b000000000000000100010010;
		16'b1110101001100001 : data_out =  24'b000000000000000100010010;
		16'b1110101001100011 : data_out =  24'b000000000000000100010010;
		16'b1110101001100101 : data_out =  24'b000000000000000100010010;
		16'b1110101001100111 : data_out =  24'b000000000000000100010011;
		16'b1110101001101001 : data_out =  24'b000000000000000100010011;
		16'b1110101001101011 : data_out =  24'b000000000000000100010011;
		16'b1110101001101101 : data_out =  24'b000000000000000100010100;
		16'b1110101001101111 : data_out =  24'b000000000000000100010100;
		16'b1110101001110001 : data_out =  24'b000000000000000100010100;
		16'b1110101001110011 : data_out =  24'b000000000000000100010100;
		16'b1110101001110101 : data_out =  24'b000000000000000100010101;
		16'b1110101001110111 : data_out =  24'b000000000000000100010101;
		16'b1110101001111001 : data_out =  24'b000000000000000100010101;
		16'b1110101001111011 : data_out =  24'b000000000000000100010110;
		16'b1110101001111101 : data_out =  24'b000000000000000100010110;
		16'b1110101001111111 : data_out =  24'b000000000000000100010110;
		16'b1110101010000010 : data_out =  24'b000000000000000100010110;
		16'b1110101010000100 : data_out =  24'b000000000000000100010111;
		16'b1110101010000110 : data_out =  24'b000000000000000100010111;
		16'b1110101010001000 : data_out =  24'b000000000000000100010111;
		16'b1110101010001010 : data_out =  24'b000000000000000100010111;
		16'b1110101010001100 : data_out =  24'b000000000000000100011000;
		16'b1110101010001110 : data_out =  24'b000000000000000100011000;
		16'b1110101010010000 : data_out =  24'b000000000000000100011000;
		16'b1110101010010010 : data_out =  24'b000000000000000100011001;
		16'b1110101010010100 : data_out =  24'b000000000000000100011001;
		16'b1110101010010110 : data_out =  24'b000000000000000100011001;
		16'b1110101010011000 : data_out =  24'b000000000000000100011001;
		16'b1110101010011010 : data_out =  24'b000000000000000100011010;
		16'b1110101010011100 : data_out =  24'b000000000000000100011010;
		16'b1110101010011110 : data_out =  24'b000000000000000100011010;
		16'b1110101010100000 : data_out =  24'b000000000000000100011011;
		16'b1110101010100010 : data_out =  24'b000000000000000100011011;
		16'b1110101010100100 : data_out =  24'b000000000000000100011011;
		16'b1110101010100110 : data_out =  24'b000000000000000100011011;
		16'b1110101010101000 : data_out =  24'b000000000000000100011100;
		16'b1110101010101010 : data_out =  24'b000000000000000100011100;
		16'b1110101010101101 : data_out =  24'b000000000000000100011100;
		16'b1110101010101111 : data_out =  24'b000000000000000100011101;
		16'b1110101010110001 : data_out =  24'b000000000000000100011101;
		16'b1110101010110011 : data_out =  24'b000000000000000100011101;
		16'b1110101010110101 : data_out =  24'b000000000000000100011101;
		16'b1110101010110111 : data_out =  24'b000000000000000100011110;
		16'b1110101010111001 : data_out =  24'b000000000000000100011110;
		16'b1110101010111011 : data_out =  24'b000000000000000100011110;
		16'b1110101010111101 : data_out =  24'b000000000000000100011111;
		16'b1110101010111111 : data_out =  24'b000000000000000100011111;
		16'b1110101011000001 : data_out =  24'b000000000000000100011111;
		16'b1110101011000011 : data_out =  24'b000000000000000100011111;
		16'b1110101011000101 : data_out =  24'b000000000000000100100000;
		16'b1110101011000111 : data_out =  24'b000000000000000100100000;
		16'b1110101011001001 : data_out =  24'b000000000000000100100000;
		16'b1110101011001011 : data_out =  24'b000000000000000100100001;
		16'b1110101011001101 : data_out =  24'b000000000000000100100001;
		16'b1110101011001111 : data_out =  24'b000000000000000100100001;
		16'b1110101011010001 : data_out =  24'b000000000000000100100001;
		16'b1110101011010011 : data_out =  24'b000000000000000100100010;
		16'b1110101011010101 : data_out =  24'b000000000000000100100010;
		16'b1110101011011000 : data_out =  24'b000000000000000100100010;
		16'b1110101011011010 : data_out =  24'b000000000000000100100011;
		16'b1110101011011100 : data_out =  24'b000000000000000100100011;
		16'b1110101011011110 : data_out =  24'b000000000000000100100011;
		16'b1110101011100000 : data_out =  24'b000000000000000100100100;
		16'b1110101011100010 : data_out =  24'b000000000000000100100100;
		16'b1110101011100100 : data_out =  24'b000000000000000100100100;
		16'b1110101011100110 : data_out =  24'b000000000000000100100100;
		16'b1110101011101000 : data_out =  24'b000000000000000100100101;
		16'b1110101011101010 : data_out =  24'b000000000000000100100101;
		16'b1110101011101100 : data_out =  24'b000000000000000100100101;
		16'b1110101011101110 : data_out =  24'b000000000000000100100110;
		16'b1110101011110000 : data_out =  24'b000000000000000100100110;
		16'b1110101011110010 : data_out =  24'b000000000000000100100110;
		16'b1110101011110100 : data_out =  24'b000000000000000100100110;
		16'b1110101011110110 : data_out =  24'b000000000000000100100111;
		16'b1110101011111000 : data_out =  24'b000000000000000100100111;
		16'b1110101011111010 : data_out =  24'b000000000000000100100111;
		16'b1110101011111100 : data_out =  24'b000000000000000100101000;
		16'b1110101011111110 : data_out =  24'b000000000000000100101000;
		16'b1110101100000001 : data_out =  24'b000000000000000100101000;
		16'b1110101100000011 : data_out =  24'b000000000000000100101001;
		16'b1110101100000101 : data_out =  24'b000000000000000100101001;
		16'b1110101100000111 : data_out =  24'b000000000000000100101001;
		16'b1110101100001001 : data_out =  24'b000000000000000100101001;
		16'b1110101100001011 : data_out =  24'b000000000000000100101010;
		16'b1110101100001101 : data_out =  24'b000000000000000100101010;
		16'b1110101100001111 : data_out =  24'b000000000000000100101010;
		16'b1110101100010001 : data_out =  24'b000000000000000100101011;
		16'b1110101100010011 : data_out =  24'b000000000000000100101011;
		16'b1110101100010101 : data_out =  24'b000000000000000100101011;
		16'b1110101100010111 : data_out =  24'b000000000000000100101011;
		16'b1110101100011001 : data_out =  24'b000000000000000100101100;
		16'b1110101100011011 : data_out =  24'b000000000000000100101100;
		16'b1110101100011101 : data_out =  24'b000000000000000100101100;
		16'b1110101100011111 : data_out =  24'b000000000000000100101101;
		16'b1110101100100001 : data_out =  24'b000000000000000100101101;
		16'b1110101100100011 : data_out =  24'b000000000000000100101101;
		16'b1110101100100101 : data_out =  24'b000000000000000100101110;
		16'b1110101100100111 : data_out =  24'b000000000000000100101110;
		16'b1110101100101001 : data_out =  24'b000000000000000100101110;
		16'b1110101100101100 : data_out =  24'b000000000000000100101111;
		16'b1110101100101110 : data_out =  24'b000000000000000100101111;
		16'b1110101100110000 : data_out =  24'b000000000000000100101111;
		16'b1110101100110010 : data_out =  24'b000000000000000100101111;
		16'b1110101100110100 : data_out =  24'b000000000000000100110000;
		16'b1110101100110110 : data_out =  24'b000000000000000100110000;
		16'b1110101100111000 : data_out =  24'b000000000000000100110000;
		16'b1110101100111010 : data_out =  24'b000000000000000100110001;
		16'b1110101100111100 : data_out =  24'b000000000000000100110001;
		16'b1110101100111110 : data_out =  24'b000000000000000100110001;
		16'b1110101101000000 : data_out =  24'b000000000000000100110010;
		16'b1110101101000010 : data_out =  24'b000000000000000100110010;
		16'b1110101101000100 : data_out =  24'b000000000000000100110010;
		16'b1110101101000110 : data_out =  24'b000000000000000100110010;
		16'b1110101101001000 : data_out =  24'b000000000000000100110011;
		16'b1110101101001010 : data_out =  24'b000000000000000100110011;
		16'b1110101101001100 : data_out =  24'b000000000000000100110011;
		16'b1110101101001110 : data_out =  24'b000000000000000100110100;
		16'b1110101101010000 : data_out =  24'b000000000000000100110100;
		16'b1110101101010010 : data_out =  24'b000000000000000100110100;
		16'b1110101101010100 : data_out =  24'b000000000000000100110101;
		16'b1110101101010111 : data_out =  24'b000000000000000100110101;
		16'b1110101101011001 : data_out =  24'b000000000000000100110101;
		16'b1110101101011011 : data_out =  24'b000000000000000100110110;
		16'b1110101101011101 : data_out =  24'b000000000000000100110110;
		16'b1110101101011111 : data_out =  24'b000000000000000100110110;
		16'b1110101101100001 : data_out =  24'b000000000000000100110110;
		16'b1110101101100011 : data_out =  24'b000000000000000100110111;
		16'b1110101101100101 : data_out =  24'b000000000000000100110111;
		16'b1110101101100111 : data_out =  24'b000000000000000100110111;
		16'b1110101101101001 : data_out =  24'b000000000000000100111000;
		16'b1110101101101011 : data_out =  24'b000000000000000100111000;
		16'b1110101101101101 : data_out =  24'b000000000000000100111000;
		16'b1110101101101111 : data_out =  24'b000000000000000100111001;
		16'b1110101101110001 : data_out =  24'b000000000000000100111001;
		16'b1110101101110011 : data_out =  24'b000000000000000100111001;
		16'b1110101101110101 : data_out =  24'b000000000000000100111010;
		16'b1110101101110111 : data_out =  24'b000000000000000100111010;
		16'b1110101101111001 : data_out =  24'b000000000000000100111010;
		16'b1110101101111011 : data_out =  24'b000000000000000100111011;
		16'b1110101101111101 : data_out =  24'b000000000000000100111011;
		16'b1110101101111111 : data_out =  24'b000000000000000100111011;
		16'b1110101110000010 : data_out =  24'b000000000000000100111100;
		16'b1110101110000100 : data_out =  24'b000000000000000100111100;
		16'b1110101110000110 : data_out =  24'b000000000000000100111100;
		16'b1110101110001000 : data_out =  24'b000000000000000100111100;
		16'b1110101110001010 : data_out =  24'b000000000000000100111101;
		16'b1110101110001100 : data_out =  24'b000000000000000100111101;
		16'b1110101110001110 : data_out =  24'b000000000000000100111101;
		16'b1110101110010000 : data_out =  24'b000000000000000100111110;
		16'b1110101110010010 : data_out =  24'b000000000000000100111110;
		16'b1110101110010100 : data_out =  24'b000000000000000100111110;
		16'b1110101110010110 : data_out =  24'b000000000000000100111111;
		16'b1110101110011000 : data_out =  24'b000000000000000100111111;
		16'b1110101110011010 : data_out =  24'b000000000000000100111111;
		16'b1110101110011100 : data_out =  24'b000000000000000101000000;
		16'b1110101110011110 : data_out =  24'b000000000000000101000000;
		16'b1110101110100000 : data_out =  24'b000000000000000101000000;
		16'b1110101110100010 : data_out =  24'b000000000000000101000001;
		16'b1110101110100100 : data_out =  24'b000000000000000101000001;
		16'b1110101110100110 : data_out =  24'b000000000000000101000001;
		16'b1110101110101000 : data_out =  24'b000000000000000101000010;
		16'b1110101110101010 : data_out =  24'b000000000000000101000010;
		16'b1110101110101101 : data_out =  24'b000000000000000101000010;
		16'b1110101110101111 : data_out =  24'b000000000000000101000011;
		16'b1110101110110001 : data_out =  24'b000000000000000101000011;
		16'b1110101110110011 : data_out =  24'b000000000000000101000011;
		16'b1110101110110101 : data_out =  24'b000000000000000101000100;
		16'b1110101110110111 : data_out =  24'b000000000000000101000100;
		16'b1110101110111001 : data_out =  24'b000000000000000101000100;
		16'b1110101110111011 : data_out =  24'b000000000000000101000100;
		16'b1110101110111101 : data_out =  24'b000000000000000101000101;
		16'b1110101110111111 : data_out =  24'b000000000000000101000101;
		16'b1110101111000001 : data_out =  24'b000000000000000101000101;
		16'b1110101111000011 : data_out =  24'b000000000000000101000110;
		16'b1110101111000101 : data_out =  24'b000000000000000101000110;
		16'b1110101111000111 : data_out =  24'b000000000000000101000110;
		16'b1110101111001001 : data_out =  24'b000000000000000101000111;
		16'b1110101111001011 : data_out =  24'b000000000000000101000111;
		16'b1110101111001101 : data_out =  24'b000000000000000101000111;
		16'b1110101111001111 : data_out =  24'b000000000000000101001000;
		16'b1110101111010001 : data_out =  24'b000000000000000101001000;
		16'b1110101111010011 : data_out =  24'b000000000000000101001000;
		16'b1110101111010101 : data_out =  24'b000000000000000101001001;
		16'b1110101111011000 : data_out =  24'b000000000000000101001001;
		16'b1110101111011010 : data_out =  24'b000000000000000101001001;
		16'b1110101111011100 : data_out =  24'b000000000000000101001010;
		16'b1110101111011110 : data_out =  24'b000000000000000101001010;
		16'b1110101111100000 : data_out =  24'b000000000000000101001010;
		16'b1110101111100010 : data_out =  24'b000000000000000101001011;
		16'b1110101111100100 : data_out =  24'b000000000000000101001011;
		16'b1110101111100110 : data_out =  24'b000000000000000101001011;
		16'b1110101111101000 : data_out =  24'b000000000000000101001100;
		16'b1110101111101010 : data_out =  24'b000000000000000101001100;
		16'b1110101111101100 : data_out =  24'b000000000000000101001100;
		16'b1110101111101110 : data_out =  24'b000000000000000101001101;
		16'b1110101111110000 : data_out =  24'b000000000000000101001101;
		16'b1110101111110010 : data_out =  24'b000000000000000101001101;
		16'b1110101111110100 : data_out =  24'b000000000000000101001110;
		16'b1110101111110110 : data_out =  24'b000000000000000101001110;
		16'b1110101111111000 : data_out =  24'b000000000000000101001110;
		16'b1110101111111010 : data_out =  24'b000000000000000101001111;
		16'b1110101111111100 : data_out =  24'b000000000000000101001111;
		16'b1110101111111110 : data_out =  24'b000000000000000101001111;
		16'b1110110000000001 : data_out =  24'b000000000000000101010000;
		16'b1110110000000011 : data_out =  24'b000000000000000101010000;
		16'b1110110000000101 : data_out =  24'b000000000000000101010000;
		16'b1110110000000111 : data_out =  24'b000000000000000101010001;
		16'b1110110000001001 : data_out =  24'b000000000000000101010001;
		16'b1110110000001011 : data_out =  24'b000000000000000101010001;
		16'b1110110000001101 : data_out =  24'b000000000000000101010010;
		16'b1110110000001111 : data_out =  24'b000000000000000101010010;
		16'b1110110000010001 : data_out =  24'b000000000000000101010010;
		16'b1110110000010011 : data_out =  24'b000000000000000101010011;
		16'b1110110000010101 : data_out =  24'b000000000000000101010011;
		16'b1110110000010111 : data_out =  24'b000000000000000101010011;
		16'b1110110000011001 : data_out =  24'b000000000000000101010100;
		16'b1110110000011011 : data_out =  24'b000000000000000101010100;
		16'b1110110000011101 : data_out =  24'b000000000000000101010100;
		16'b1110110000011111 : data_out =  24'b000000000000000101010101;
		16'b1110110000100001 : data_out =  24'b000000000000000101010101;
		16'b1110110000100011 : data_out =  24'b000000000000000101010101;
		16'b1110110000100101 : data_out =  24'b000000000000000101010110;
		16'b1110110000100111 : data_out =  24'b000000000000000101010110;
		16'b1110110000101001 : data_out =  24'b000000000000000101010111;
		16'b1110110000101100 : data_out =  24'b000000000000000101010111;
		16'b1110110000101110 : data_out =  24'b000000000000000101010111;
		16'b1110110000110000 : data_out =  24'b000000000000000101011000;
		16'b1110110000110010 : data_out =  24'b000000000000000101011000;
		16'b1110110000110100 : data_out =  24'b000000000000000101011000;
		16'b1110110000110110 : data_out =  24'b000000000000000101011001;
		16'b1110110000111000 : data_out =  24'b000000000000000101011001;
		16'b1110110000111010 : data_out =  24'b000000000000000101011001;
		16'b1110110000111100 : data_out =  24'b000000000000000101011010;
		16'b1110110000111110 : data_out =  24'b000000000000000101011010;
		16'b1110110001000000 : data_out =  24'b000000000000000101011010;
		16'b1110110001000010 : data_out =  24'b000000000000000101011011;
		16'b1110110001000100 : data_out =  24'b000000000000000101011011;
		16'b1110110001000110 : data_out =  24'b000000000000000101011011;
		16'b1110110001001000 : data_out =  24'b000000000000000101011100;
		16'b1110110001001010 : data_out =  24'b000000000000000101011100;
		16'b1110110001001100 : data_out =  24'b000000000000000101011100;
		16'b1110110001001110 : data_out =  24'b000000000000000101011101;
		16'b1110110001010000 : data_out =  24'b000000000000000101011101;
		16'b1110110001010010 : data_out =  24'b000000000000000101011101;
		16'b1110110001010100 : data_out =  24'b000000000000000101011110;
		16'b1110110001010111 : data_out =  24'b000000000000000101011110;
		16'b1110110001011001 : data_out =  24'b000000000000000101011110;
		16'b1110110001011011 : data_out =  24'b000000000000000101011111;
		16'b1110110001011101 : data_out =  24'b000000000000000101011111;
		16'b1110110001011111 : data_out =  24'b000000000000000101100000;
		16'b1110110001100001 : data_out =  24'b000000000000000101100000;
		16'b1110110001100011 : data_out =  24'b000000000000000101100000;
		16'b1110110001100101 : data_out =  24'b000000000000000101100001;
		16'b1110110001100111 : data_out =  24'b000000000000000101100001;
		16'b1110110001101001 : data_out =  24'b000000000000000101100001;
		16'b1110110001101011 : data_out =  24'b000000000000000101100010;
		16'b1110110001101101 : data_out =  24'b000000000000000101100010;
		16'b1110110001101111 : data_out =  24'b000000000000000101100010;
		16'b1110110001110001 : data_out =  24'b000000000000000101100011;
		16'b1110110001110011 : data_out =  24'b000000000000000101100011;
		16'b1110110001110101 : data_out =  24'b000000000000000101100011;
		16'b1110110001110111 : data_out =  24'b000000000000000101100100;
		16'b1110110001111001 : data_out =  24'b000000000000000101100100;
		16'b1110110001111011 : data_out =  24'b000000000000000101100101;
		16'b1110110001111101 : data_out =  24'b000000000000000101100101;
		16'b1110110001111111 : data_out =  24'b000000000000000101100101;
		16'b1110110010000010 : data_out =  24'b000000000000000101100110;
		16'b1110110010000100 : data_out =  24'b000000000000000101100110;
		16'b1110110010000110 : data_out =  24'b000000000000000101100110;
		16'b1110110010001000 : data_out =  24'b000000000000000101100111;
		16'b1110110010001010 : data_out =  24'b000000000000000101100111;
		16'b1110110010001100 : data_out =  24'b000000000000000101100111;
		16'b1110110010001110 : data_out =  24'b000000000000000101101000;
		16'b1110110010010000 : data_out =  24'b000000000000000101101000;
		16'b1110110010010010 : data_out =  24'b000000000000000101101000;
		16'b1110110010010100 : data_out =  24'b000000000000000101101001;
		16'b1110110010010110 : data_out =  24'b000000000000000101101001;
		16'b1110110010011000 : data_out =  24'b000000000000000101101010;
		16'b1110110010011010 : data_out =  24'b000000000000000101101010;
		16'b1110110010011100 : data_out =  24'b000000000000000101101010;
		16'b1110110010011110 : data_out =  24'b000000000000000101101011;
		16'b1110110010100000 : data_out =  24'b000000000000000101101011;
		16'b1110110010100010 : data_out =  24'b000000000000000101101011;
		16'b1110110010100100 : data_out =  24'b000000000000000101101100;
		16'b1110110010100110 : data_out =  24'b000000000000000101101100;
		16'b1110110010101000 : data_out =  24'b000000000000000101101100;
		16'b1110110010101010 : data_out =  24'b000000000000000101101101;
		16'b1110110010101101 : data_out =  24'b000000000000000101101101;
		16'b1110110010101111 : data_out =  24'b000000000000000101101110;
		16'b1110110010110001 : data_out =  24'b000000000000000101101110;
		16'b1110110010110011 : data_out =  24'b000000000000000101101110;
		16'b1110110010110101 : data_out =  24'b000000000000000101101111;
		16'b1110110010110111 : data_out =  24'b000000000000000101101111;
		16'b1110110010111001 : data_out =  24'b000000000000000101101111;
		16'b1110110010111011 : data_out =  24'b000000000000000101110000;
		16'b1110110010111101 : data_out =  24'b000000000000000101110000;
		16'b1110110010111111 : data_out =  24'b000000000000000101110000;
		16'b1110110011000001 : data_out =  24'b000000000000000101110001;
		16'b1110110011000011 : data_out =  24'b000000000000000101110001;
		16'b1110110011000101 : data_out =  24'b000000000000000101110010;
		16'b1110110011000111 : data_out =  24'b000000000000000101110010;
		16'b1110110011001001 : data_out =  24'b000000000000000101110010;
		16'b1110110011001011 : data_out =  24'b000000000000000101110011;
		16'b1110110011001101 : data_out =  24'b000000000000000101110011;
		16'b1110110011001111 : data_out =  24'b000000000000000101110011;
		16'b1110110011010001 : data_out =  24'b000000000000000101110100;
		16'b1110110011010011 : data_out =  24'b000000000000000101110100;
		16'b1110110011010101 : data_out =  24'b000000000000000101110101;
		16'b1110110011011000 : data_out =  24'b000000000000000101110101;
		16'b1110110011011010 : data_out =  24'b000000000000000101110101;
		16'b1110110011011100 : data_out =  24'b000000000000000101110110;
		16'b1110110011011110 : data_out =  24'b000000000000000101110110;
		16'b1110110011100000 : data_out =  24'b000000000000000101110110;
		16'b1110110011100010 : data_out =  24'b000000000000000101110111;
		16'b1110110011100100 : data_out =  24'b000000000000000101110111;
		16'b1110110011100110 : data_out =  24'b000000000000000101111000;
		16'b1110110011101000 : data_out =  24'b000000000000000101111000;
		16'b1110110011101010 : data_out =  24'b000000000000000101111000;
		16'b1110110011101100 : data_out =  24'b000000000000000101111001;
		16'b1110110011101110 : data_out =  24'b000000000000000101111001;
		16'b1110110011110000 : data_out =  24'b000000000000000101111001;
		16'b1110110011110010 : data_out =  24'b000000000000000101111010;
		16'b1110110011110100 : data_out =  24'b000000000000000101111010;
		16'b1110110011110110 : data_out =  24'b000000000000000101111011;
		16'b1110110011111000 : data_out =  24'b000000000000000101111011;
		16'b1110110011111010 : data_out =  24'b000000000000000101111011;
		16'b1110110011111100 : data_out =  24'b000000000000000101111100;
		16'b1110110011111110 : data_out =  24'b000000000000000101111100;
		16'b1110110100000001 : data_out =  24'b000000000000000101111100;
		16'b1110110100000011 : data_out =  24'b000000000000000101111101;
		16'b1110110100000101 : data_out =  24'b000000000000000101111101;
		16'b1110110100000111 : data_out =  24'b000000000000000101111110;
		16'b1110110100001001 : data_out =  24'b000000000000000101111110;
		16'b1110110100001011 : data_out =  24'b000000000000000101111110;
		16'b1110110100001101 : data_out =  24'b000000000000000101111111;
		16'b1110110100001111 : data_out =  24'b000000000000000101111111;
		16'b1110110100010001 : data_out =  24'b000000000000000110000000;
		16'b1110110100010011 : data_out =  24'b000000000000000110000000;
		16'b1110110100010101 : data_out =  24'b000000000000000110000000;
		16'b1110110100010111 : data_out =  24'b000000000000000110000001;
		16'b1110110100011001 : data_out =  24'b000000000000000110000001;
		16'b1110110100011011 : data_out =  24'b000000000000000110000001;
		16'b1110110100011101 : data_out =  24'b000000000000000110000010;
		16'b1110110100011111 : data_out =  24'b000000000000000110000010;
		16'b1110110100100001 : data_out =  24'b000000000000000110000011;
		16'b1110110100100011 : data_out =  24'b000000000000000110000011;
		16'b1110110100100101 : data_out =  24'b000000000000000110000011;
		16'b1110110100100111 : data_out =  24'b000000000000000110000100;
		16'b1110110100101001 : data_out =  24'b000000000000000110000100;
		16'b1110110100101100 : data_out =  24'b000000000000000110000101;
		16'b1110110100101110 : data_out =  24'b000000000000000110000101;
		16'b1110110100110000 : data_out =  24'b000000000000000110000101;
		16'b1110110100110010 : data_out =  24'b000000000000000110000110;
		16'b1110110100110100 : data_out =  24'b000000000000000110000110;
		16'b1110110100110110 : data_out =  24'b000000000000000110000111;
		16'b1110110100111000 : data_out =  24'b000000000000000110000111;
		16'b1110110100111010 : data_out =  24'b000000000000000110000111;
		16'b1110110100111100 : data_out =  24'b000000000000000110001000;
		16'b1110110100111110 : data_out =  24'b000000000000000110001000;
		16'b1110110101000000 : data_out =  24'b000000000000000110001000;
		16'b1110110101000010 : data_out =  24'b000000000000000110001001;
		16'b1110110101000100 : data_out =  24'b000000000000000110001001;
		16'b1110110101000110 : data_out =  24'b000000000000000110001010;
		16'b1110110101001000 : data_out =  24'b000000000000000110001010;
		16'b1110110101001010 : data_out =  24'b000000000000000110001010;
		16'b1110110101001100 : data_out =  24'b000000000000000110001011;
		16'b1110110101001110 : data_out =  24'b000000000000000110001011;
		16'b1110110101010000 : data_out =  24'b000000000000000110001100;
		16'b1110110101010010 : data_out =  24'b000000000000000110001100;
		16'b1110110101010100 : data_out =  24'b000000000000000110001100;
		16'b1110110101010111 : data_out =  24'b000000000000000110001101;
		16'b1110110101011001 : data_out =  24'b000000000000000110001101;
		16'b1110110101011011 : data_out =  24'b000000000000000110001110;
		16'b1110110101011101 : data_out =  24'b000000000000000110001110;
		16'b1110110101011111 : data_out =  24'b000000000000000110001110;
		16'b1110110101100001 : data_out =  24'b000000000000000110001111;
		16'b1110110101100011 : data_out =  24'b000000000000000110001111;
		16'b1110110101100101 : data_out =  24'b000000000000000110010000;
		16'b1110110101100111 : data_out =  24'b000000000000000110010000;
		16'b1110110101101001 : data_out =  24'b000000000000000110010000;
		16'b1110110101101011 : data_out =  24'b000000000000000110010001;
		16'b1110110101101101 : data_out =  24'b000000000000000110010001;
		16'b1110110101101111 : data_out =  24'b000000000000000110010010;
		16'b1110110101110001 : data_out =  24'b000000000000000110010010;
		16'b1110110101110011 : data_out =  24'b000000000000000110010010;
		16'b1110110101110101 : data_out =  24'b000000000000000110010011;
		16'b1110110101110111 : data_out =  24'b000000000000000110010011;
		16'b1110110101111001 : data_out =  24'b000000000000000110010100;
		16'b1110110101111011 : data_out =  24'b000000000000000110010100;
		16'b1110110101111101 : data_out =  24'b000000000000000110010100;
		16'b1110110101111111 : data_out =  24'b000000000000000110010101;
		16'b1110110110000010 : data_out =  24'b000000000000000110010101;
		16'b1110110110000100 : data_out =  24'b000000000000000110010110;
		16'b1110110110000110 : data_out =  24'b000000000000000110010110;
		16'b1110110110001000 : data_out =  24'b000000000000000110010110;
		16'b1110110110001010 : data_out =  24'b000000000000000110010111;
		16'b1110110110001100 : data_out =  24'b000000000000000110010111;
		16'b1110110110001110 : data_out =  24'b000000000000000110011000;
		16'b1110110110010000 : data_out =  24'b000000000000000110011000;
		16'b1110110110010010 : data_out =  24'b000000000000000110011001;
		16'b1110110110010100 : data_out =  24'b000000000000000110011001;
		16'b1110110110010110 : data_out =  24'b000000000000000110011001;
		16'b1110110110011000 : data_out =  24'b000000000000000110011010;
		16'b1110110110011010 : data_out =  24'b000000000000000110011010;
		16'b1110110110011100 : data_out =  24'b000000000000000110011011;
		16'b1110110110011110 : data_out =  24'b000000000000000110011011;
		16'b1110110110100000 : data_out =  24'b000000000000000110011011;
		16'b1110110110100010 : data_out =  24'b000000000000000110011100;
		16'b1110110110100100 : data_out =  24'b000000000000000110011100;
		16'b1110110110100110 : data_out =  24'b000000000000000110011101;
		16'b1110110110101000 : data_out =  24'b000000000000000110011101;
		16'b1110110110101010 : data_out =  24'b000000000000000110011101;
		16'b1110110110101101 : data_out =  24'b000000000000000110011110;
		16'b1110110110101111 : data_out =  24'b000000000000000110011110;
		16'b1110110110110001 : data_out =  24'b000000000000000110011111;
		16'b1110110110110011 : data_out =  24'b000000000000000110011111;
		16'b1110110110110101 : data_out =  24'b000000000000000110100000;
		16'b1110110110110111 : data_out =  24'b000000000000000110100000;
		16'b1110110110111001 : data_out =  24'b000000000000000110100000;
		16'b1110110110111011 : data_out =  24'b000000000000000110100001;
		16'b1110110110111101 : data_out =  24'b000000000000000110100001;
		16'b1110110110111111 : data_out =  24'b000000000000000110100010;
		16'b1110110111000001 : data_out =  24'b000000000000000110100010;
		16'b1110110111000011 : data_out =  24'b000000000000000110100010;
		16'b1110110111000101 : data_out =  24'b000000000000000110100011;
		16'b1110110111000111 : data_out =  24'b000000000000000110100011;
		16'b1110110111001001 : data_out =  24'b000000000000000110100100;
		16'b1110110111001011 : data_out =  24'b000000000000000110100100;
		16'b1110110111001101 : data_out =  24'b000000000000000110100101;
		16'b1110110111001111 : data_out =  24'b000000000000000110100101;
		16'b1110110111010001 : data_out =  24'b000000000000000110100101;
		16'b1110110111010011 : data_out =  24'b000000000000000110100110;
		16'b1110110111010101 : data_out =  24'b000000000000000110100110;
		16'b1110110111011000 : data_out =  24'b000000000000000110100111;
		16'b1110110111011010 : data_out =  24'b000000000000000110100111;
		16'b1110110111011100 : data_out =  24'b000000000000000110101000;
		16'b1110110111011110 : data_out =  24'b000000000000000110101000;
		16'b1110110111100000 : data_out =  24'b000000000000000110101000;
		16'b1110110111100010 : data_out =  24'b000000000000000110101001;
		16'b1110110111100100 : data_out =  24'b000000000000000110101001;
		16'b1110110111100110 : data_out =  24'b000000000000000110101010;
		16'b1110110111101000 : data_out =  24'b000000000000000110101010;
		16'b1110110111101010 : data_out =  24'b000000000000000110101010;
		16'b1110110111101100 : data_out =  24'b000000000000000110101011;
		16'b1110110111101110 : data_out =  24'b000000000000000110101011;
		16'b1110110111110000 : data_out =  24'b000000000000000110101100;
		16'b1110110111110010 : data_out =  24'b000000000000000110101100;
		16'b1110110111110100 : data_out =  24'b000000000000000110101101;
		16'b1110110111110110 : data_out =  24'b000000000000000110101101;
		16'b1110110111111000 : data_out =  24'b000000000000000110101101;
		16'b1110110111111010 : data_out =  24'b000000000000000110101110;
		16'b1110110111111100 : data_out =  24'b000000000000000110101110;
		16'b1110110111111110 : data_out =  24'b000000000000000110101111;
		16'b1110111000000001 : data_out =  24'b000000000000000110101111;
		16'b1110111000000011 : data_out =  24'b000000000000000110110000;
		16'b1110111000000101 : data_out =  24'b000000000000000110110000;
		16'b1110111000000111 : data_out =  24'b000000000000000110110001;
		16'b1110111000001001 : data_out =  24'b000000000000000110110001;
		16'b1110111000001011 : data_out =  24'b000000000000000110110001;
		16'b1110111000001101 : data_out =  24'b000000000000000110110010;
		16'b1110111000001111 : data_out =  24'b000000000000000110110010;
		16'b1110111000010001 : data_out =  24'b000000000000000110110011;
		16'b1110111000010011 : data_out =  24'b000000000000000110110011;
		16'b1110111000010101 : data_out =  24'b000000000000000110110100;
		16'b1110111000010111 : data_out =  24'b000000000000000110110100;
		16'b1110111000011001 : data_out =  24'b000000000000000110110100;
		16'b1110111000011011 : data_out =  24'b000000000000000110110101;
		16'b1110111000011101 : data_out =  24'b000000000000000110110101;
		16'b1110111000011111 : data_out =  24'b000000000000000110110110;
		16'b1110111000100001 : data_out =  24'b000000000000000110110110;
		16'b1110111000100011 : data_out =  24'b000000000000000110110111;
		16'b1110111000100101 : data_out =  24'b000000000000000110110111;
		16'b1110111000100111 : data_out =  24'b000000000000000110110111;
		16'b1110111000101001 : data_out =  24'b000000000000000110111000;
		16'b1110111000101100 : data_out =  24'b000000000000000110111000;
		16'b1110111000101110 : data_out =  24'b000000000000000110111001;
		16'b1110111000110000 : data_out =  24'b000000000000000110111001;
		16'b1110111000110010 : data_out =  24'b000000000000000110111010;
		16'b1110111000110100 : data_out =  24'b000000000000000110111010;
		16'b1110111000110110 : data_out =  24'b000000000000000110111011;
		16'b1110111000111000 : data_out =  24'b000000000000000110111011;
		16'b1110111000111010 : data_out =  24'b000000000000000110111011;
		16'b1110111000111100 : data_out =  24'b000000000000000110111100;
		16'b1110111000111110 : data_out =  24'b000000000000000110111100;
		16'b1110111001000000 : data_out =  24'b000000000000000110111101;
		16'b1110111001000010 : data_out =  24'b000000000000000110111101;
		16'b1110111001000100 : data_out =  24'b000000000000000110111110;
		16'b1110111001000110 : data_out =  24'b000000000000000110111110;
		16'b1110111001001000 : data_out =  24'b000000000000000110111111;
		16'b1110111001001010 : data_out =  24'b000000000000000110111111;
		16'b1110111001001100 : data_out =  24'b000000000000000110111111;
		16'b1110111001001110 : data_out =  24'b000000000000000111000000;
		16'b1110111001010000 : data_out =  24'b000000000000000111000000;
		16'b1110111001010010 : data_out =  24'b000000000000000111000001;
		16'b1110111001010100 : data_out =  24'b000000000000000111000001;
		16'b1110111001010111 : data_out =  24'b000000000000000111000010;
		16'b1110111001011001 : data_out =  24'b000000000000000111000010;
		16'b1110111001011011 : data_out =  24'b000000000000000111000011;
		16'b1110111001011101 : data_out =  24'b000000000000000111000011;
		16'b1110111001011111 : data_out =  24'b000000000000000111000100;
		16'b1110111001100001 : data_out =  24'b000000000000000111000100;
		16'b1110111001100011 : data_out =  24'b000000000000000111000100;
		16'b1110111001100101 : data_out =  24'b000000000000000111000101;
		16'b1110111001100111 : data_out =  24'b000000000000000111000101;
		16'b1110111001101001 : data_out =  24'b000000000000000111000110;
		16'b1110111001101011 : data_out =  24'b000000000000000111000110;
		16'b1110111001101101 : data_out =  24'b000000000000000111000111;
		16'b1110111001101111 : data_out =  24'b000000000000000111000111;
		16'b1110111001110001 : data_out =  24'b000000000000000111001000;
		16'b1110111001110011 : data_out =  24'b000000000000000111001000;
		16'b1110111001110101 : data_out =  24'b000000000000000111001001;
		16'b1110111001110111 : data_out =  24'b000000000000000111001001;
		16'b1110111001111001 : data_out =  24'b000000000000000111001001;
		16'b1110111001111011 : data_out =  24'b000000000000000111001010;
		16'b1110111001111101 : data_out =  24'b000000000000000111001010;
		16'b1110111001111111 : data_out =  24'b000000000000000111001011;
		16'b1110111010000010 : data_out =  24'b000000000000000111001011;
		16'b1110111010000100 : data_out =  24'b000000000000000111001100;
		16'b1110111010000110 : data_out =  24'b000000000000000111001100;
		16'b1110111010001000 : data_out =  24'b000000000000000111001101;
		16'b1110111010001010 : data_out =  24'b000000000000000111001101;
		16'b1110111010001100 : data_out =  24'b000000000000000111001110;
		16'b1110111010001110 : data_out =  24'b000000000000000111001110;
		16'b1110111010010000 : data_out =  24'b000000000000000111001111;
		16'b1110111010010010 : data_out =  24'b000000000000000111001111;
		16'b1110111010010100 : data_out =  24'b000000000000000111001111;
		16'b1110111010010110 : data_out =  24'b000000000000000111010000;
		16'b1110111010011000 : data_out =  24'b000000000000000111010000;
		16'b1110111010011010 : data_out =  24'b000000000000000111010001;
		16'b1110111010011100 : data_out =  24'b000000000000000111010001;
		16'b1110111010011110 : data_out =  24'b000000000000000111010010;
		16'b1110111010100000 : data_out =  24'b000000000000000111010010;
		16'b1110111010100010 : data_out =  24'b000000000000000111010011;
		16'b1110111010100100 : data_out =  24'b000000000000000111010011;
		16'b1110111010100110 : data_out =  24'b000000000000000111010100;
		16'b1110111010101000 : data_out =  24'b000000000000000111010100;
		16'b1110111010101010 : data_out =  24'b000000000000000111010101;
		16'b1110111010101101 : data_out =  24'b000000000000000111010101;
		16'b1110111010101111 : data_out =  24'b000000000000000111010110;
		16'b1110111010110001 : data_out =  24'b000000000000000111010110;
		16'b1110111010110011 : data_out =  24'b000000000000000111010110;
		16'b1110111010110101 : data_out =  24'b000000000000000111010111;
		16'b1110111010110111 : data_out =  24'b000000000000000111010111;
		16'b1110111010111001 : data_out =  24'b000000000000000111011000;
		16'b1110111010111011 : data_out =  24'b000000000000000111011000;
		16'b1110111010111101 : data_out =  24'b000000000000000111011001;
		16'b1110111010111111 : data_out =  24'b000000000000000111011001;
		16'b1110111011000001 : data_out =  24'b000000000000000111011010;
		16'b1110111011000011 : data_out =  24'b000000000000000111011010;
		16'b1110111011000101 : data_out =  24'b000000000000000111011011;
		16'b1110111011000111 : data_out =  24'b000000000000000111011011;
		16'b1110111011001001 : data_out =  24'b000000000000000111011100;
		16'b1110111011001011 : data_out =  24'b000000000000000111011100;
		16'b1110111011001101 : data_out =  24'b000000000000000111011101;
		16'b1110111011001111 : data_out =  24'b000000000000000111011101;
		16'b1110111011010001 : data_out =  24'b000000000000000111011110;
		16'b1110111011010011 : data_out =  24'b000000000000000111011110;
		16'b1110111011010101 : data_out =  24'b000000000000000111011111;
		16'b1110111011011000 : data_out =  24'b000000000000000111011111;
		16'b1110111011011010 : data_out =  24'b000000000000000111011111;
		16'b1110111011011100 : data_out =  24'b000000000000000111100000;
		16'b1110111011011110 : data_out =  24'b000000000000000111100000;
		16'b1110111011100000 : data_out =  24'b000000000000000111100001;
		16'b1110111011100010 : data_out =  24'b000000000000000111100001;
		16'b1110111011100100 : data_out =  24'b000000000000000111100010;
		16'b1110111011100110 : data_out =  24'b000000000000000111100010;
		16'b1110111011101000 : data_out =  24'b000000000000000111100011;
		16'b1110111011101010 : data_out =  24'b000000000000000111100011;
		16'b1110111011101100 : data_out =  24'b000000000000000111100100;
		16'b1110111011101110 : data_out =  24'b000000000000000111100100;
		16'b1110111011110000 : data_out =  24'b000000000000000111100101;
		16'b1110111011110010 : data_out =  24'b000000000000000111100101;
		16'b1110111011110100 : data_out =  24'b000000000000000111100110;
		16'b1110111011110110 : data_out =  24'b000000000000000111100110;
		16'b1110111011111000 : data_out =  24'b000000000000000111100111;
		16'b1110111011111010 : data_out =  24'b000000000000000111100111;
		16'b1110111011111100 : data_out =  24'b000000000000000111101000;
		16'b1110111011111110 : data_out =  24'b000000000000000111101000;
		16'b1110111100000001 : data_out =  24'b000000000000000111101001;
		16'b1110111100000011 : data_out =  24'b000000000000000111101001;
		16'b1110111100000101 : data_out =  24'b000000000000000111101010;
		16'b1110111100000111 : data_out =  24'b000000000000000111101010;
		16'b1110111100001001 : data_out =  24'b000000000000000111101011;
		16'b1110111100001011 : data_out =  24'b000000000000000111101011;
		16'b1110111100001101 : data_out =  24'b000000000000000111101100;
		16'b1110111100001111 : data_out =  24'b000000000000000111101100;
		16'b1110111100010001 : data_out =  24'b000000000000000111101101;
		16'b1110111100010011 : data_out =  24'b000000000000000111101101;
		16'b1110111100010101 : data_out =  24'b000000000000000111101110;
		16'b1110111100010111 : data_out =  24'b000000000000000111101110;
		16'b1110111100011001 : data_out =  24'b000000000000000111101111;
		16'b1110111100011011 : data_out =  24'b000000000000000111101111;
		16'b1110111100011101 : data_out =  24'b000000000000000111110000;
		16'b1110111100011111 : data_out =  24'b000000000000000111110000;
		16'b1110111100100001 : data_out =  24'b000000000000000111110001;
		16'b1110111100100011 : data_out =  24'b000000000000000111110001;
		16'b1110111100100101 : data_out =  24'b000000000000000111110010;
		16'b1110111100100111 : data_out =  24'b000000000000000111110010;
		16'b1110111100101001 : data_out =  24'b000000000000000111110011;
		16'b1110111100101100 : data_out =  24'b000000000000000111110011;
		16'b1110111100101110 : data_out =  24'b000000000000000111110100;
		16'b1110111100110000 : data_out =  24'b000000000000000111110100;
		16'b1110111100110010 : data_out =  24'b000000000000000111110101;
		16'b1110111100110100 : data_out =  24'b000000000000000111110101;
		16'b1110111100110110 : data_out =  24'b000000000000000111110110;
		16'b1110111100111000 : data_out =  24'b000000000000000111110110;
		16'b1110111100111010 : data_out =  24'b000000000000000111110111;
		16'b1110111100111100 : data_out =  24'b000000000000000111110111;
		16'b1110111100111110 : data_out =  24'b000000000000000111111000;
		16'b1110111101000000 : data_out =  24'b000000000000000111111000;
		16'b1110111101000010 : data_out =  24'b000000000000000111111001;
		16'b1110111101000100 : data_out =  24'b000000000000000111111001;
		16'b1110111101000110 : data_out =  24'b000000000000000111111010;
		16'b1110111101001000 : data_out =  24'b000000000000000111111010;
		16'b1110111101001010 : data_out =  24'b000000000000000111111011;
		16'b1110111101001100 : data_out =  24'b000000000000000111111011;
		16'b1110111101001110 : data_out =  24'b000000000000000111111100;
		16'b1110111101010000 : data_out =  24'b000000000000000111111100;
		16'b1110111101010010 : data_out =  24'b000000000000000111111101;
		16'b1110111101010100 : data_out =  24'b000000000000000111111101;
		16'b1110111101010111 : data_out =  24'b000000000000000111111110;
		16'b1110111101011001 : data_out =  24'b000000000000000111111110;
		16'b1110111101011011 : data_out =  24'b000000000000000111111111;
		16'b1110111101011101 : data_out =  24'b000000000000000111111111;
		16'b1110111101011111 : data_out =  24'b000000000000001000000000;
		16'b1110111101100001 : data_out =  24'b000000000000001000000000;
		16'b1110111101100011 : data_out =  24'b000000000000001000000001;
		16'b1110111101100101 : data_out =  24'b000000000000001000000001;
		16'b1110111101100111 : data_out =  24'b000000000000001000000010;
		16'b1110111101101001 : data_out =  24'b000000000000001000000010;
		16'b1110111101101011 : data_out =  24'b000000000000001000000011;
		16'b1110111101101101 : data_out =  24'b000000000000001000000011;
		16'b1110111101101111 : data_out =  24'b000000000000001000000100;
		16'b1110111101110001 : data_out =  24'b000000000000001000000100;
		16'b1110111101110011 : data_out =  24'b000000000000001000000101;
		16'b1110111101110101 : data_out =  24'b000000000000001000000101;
		16'b1110111101110111 : data_out =  24'b000000000000001000000110;
		16'b1110111101111001 : data_out =  24'b000000000000001000000110;
		16'b1110111101111011 : data_out =  24'b000000000000001000000111;
		16'b1110111101111101 : data_out =  24'b000000000000001000000111;
		16'b1110111101111111 : data_out =  24'b000000000000001000001000;
		16'b1110111110000010 : data_out =  24'b000000000000001000001001;
		16'b1110111110000100 : data_out =  24'b000000000000001000001001;
		16'b1110111110000110 : data_out =  24'b000000000000001000001010;
		16'b1110111110001000 : data_out =  24'b000000000000001000001010;
		16'b1110111110001010 : data_out =  24'b000000000000001000001011;
		16'b1110111110001100 : data_out =  24'b000000000000001000001011;
		16'b1110111110001110 : data_out =  24'b000000000000001000001100;
		16'b1110111110010000 : data_out =  24'b000000000000001000001100;
		16'b1110111110010010 : data_out =  24'b000000000000001000001101;
		16'b1110111110010100 : data_out =  24'b000000000000001000001101;
		16'b1110111110010110 : data_out =  24'b000000000000001000001110;
		16'b1110111110011000 : data_out =  24'b000000000000001000001110;
		16'b1110111110011010 : data_out =  24'b000000000000001000001111;
		16'b1110111110011100 : data_out =  24'b000000000000001000001111;
		16'b1110111110011110 : data_out =  24'b000000000000001000010000;
		16'b1110111110100000 : data_out =  24'b000000000000001000010000;
		16'b1110111110100010 : data_out =  24'b000000000000001000010001;
		16'b1110111110100100 : data_out =  24'b000000000000001000010001;
		16'b1110111110100110 : data_out =  24'b000000000000001000010010;
		16'b1110111110101000 : data_out =  24'b000000000000001000010011;
		16'b1110111110101010 : data_out =  24'b000000000000001000010011;
		16'b1110111110101101 : data_out =  24'b000000000000001000010100;
		16'b1110111110101111 : data_out =  24'b000000000000001000010100;
		16'b1110111110110001 : data_out =  24'b000000000000001000010101;
		16'b1110111110110011 : data_out =  24'b000000000000001000010101;
		16'b1110111110110101 : data_out =  24'b000000000000001000010110;
		16'b1110111110110111 : data_out =  24'b000000000000001000010110;
		16'b1110111110111001 : data_out =  24'b000000000000001000010111;
		16'b1110111110111011 : data_out =  24'b000000000000001000010111;
		16'b1110111110111101 : data_out =  24'b000000000000001000011000;
		16'b1110111110111111 : data_out =  24'b000000000000001000011000;
		16'b1110111111000001 : data_out =  24'b000000000000001000011001;
		16'b1110111111000011 : data_out =  24'b000000000000001000011001;
		16'b1110111111000101 : data_out =  24'b000000000000001000011010;
		16'b1110111111000111 : data_out =  24'b000000000000001000011011;
		16'b1110111111001001 : data_out =  24'b000000000000001000011011;
		16'b1110111111001011 : data_out =  24'b000000000000001000011100;
		16'b1110111111001101 : data_out =  24'b000000000000001000011100;
		16'b1110111111001111 : data_out =  24'b000000000000001000011101;
		16'b1110111111010001 : data_out =  24'b000000000000001000011101;
		16'b1110111111010011 : data_out =  24'b000000000000001000011110;
		16'b1110111111010101 : data_out =  24'b000000000000001000011110;
		16'b1110111111011000 : data_out =  24'b000000000000001000011111;
		16'b1110111111011010 : data_out =  24'b000000000000001000011111;
		16'b1110111111011100 : data_out =  24'b000000000000001000100000;
		16'b1110111111011110 : data_out =  24'b000000000000001000100000;
		16'b1110111111100000 : data_out =  24'b000000000000001000100001;
		16'b1110111111100010 : data_out =  24'b000000000000001000100010;
		16'b1110111111100100 : data_out =  24'b000000000000001000100010;
		16'b1110111111100110 : data_out =  24'b000000000000001000100011;
		16'b1110111111101000 : data_out =  24'b000000000000001000100011;
		16'b1110111111101010 : data_out =  24'b000000000000001000100100;
		16'b1110111111101100 : data_out =  24'b000000000000001000100100;
		16'b1110111111101110 : data_out =  24'b000000000000001000100101;
		16'b1110111111110000 : data_out =  24'b000000000000001000100101;
		16'b1110111111110010 : data_out =  24'b000000000000001000100110;
		16'b1110111111110100 : data_out =  24'b000000000000001000100111;
		16'b1110111111110110 : data_out =  24'b000000000000001000100111;
		16'b1110111111111000 : data_out =  24'b000000000000001000101000;
		16'b1110111111111010 : data_out =  24'b000000000000001000101000;
		16'b1110111111111100 : data_out =  24'b000000000000001000101001;
		16'b1110111111111110 : data_out =  24'b000000000000001000101001;
		16'b1111000000000001 : data_out =  24'b000000000000001000101010;
		16'b1111000000000011 : data_out =  24'b000000000000001000101010;
		16'b1111000000000101 : data_out =  24'b000000000000001000101011;
		16'b1111000000000111 : data_out =  24'b000000000000001000101011;
		16'b1111000000001001 : data_out =  24'b000000000000001000101100;
		16'b1111000000001011 : data_out =  24'b000000000000001000101101;
		16'b1111000000001101 : data_out =  24'b000000000000001000101101;
		16'b1111000000001111 : data_out =  24'b000000000000001000101110;
		16'b1111000000010001 : data_out =  24'b000000000000001000101110;
		16'b1111000000010011 : data_out =  24'b000000000000001000101111;
		16'b1111000000010101 : data_out =  24'b000000000000001000101111;
		16'b1111000000010111 : data_out =  24'b000000000000001000110000;
		16'b1111000000011001 : data_out =  24'b000000000000001000110001;
		16'b1111000000011011 : data_out =  24'b000000000000001000110001;
		16'b1111000000011101 : data_out =  24'b000000000000001000110010;
		16'b1111000000011111 : data_out =  24'b000000000000001000110010;
		16'b1111000000100001 : data_out =  24'b000000000000001000110011;
		16'b1111000000100011 : data_out =  24'b000000000000001000110011;
		16'b1111000000100101 : data_out =  24'b000000000000001000110100;
		16'b1111000000100111 : data_out =  24'b000000000000001000110100;
		16'b1111000000101001 : data_out =  24'b000000000000001000110101;
		16'b1111000000101100 : data_out =  24'b000000000000001000110110;
		16'b1111000000101110 : data_out =  24'b000000000000001000110110;
		16'b1111000000110000 : data_out =  24'b000000000000001000110111;
		16'b1111000000110010 : data_out =  24'b000000000000001000110111;
		16'b1111000000110100 : data_out =  24'b000000000000001000111000;
		16'b1111000000110110 : data_out =  24'b000000000000001000111000;
		16'b1111000000111000 : data_out =  24'b000000000000001000111001;
		16'b1111000000111010 : data_out =  24'b000000000000001000111010;
		16'b1111000000111100 : data_out =  24'b000000000000001000111010;
		16'b1111000000111110 : data_out =  24'b000000000000001000111011;
		16'b1111000001000000 : data_out =  24'b000000000000001000111011;
		16'b1111000001000010 : data_out =  24'b000000000000001000111100;
		16'b1111000001000100 : data_out =  24'b000000000000001000111100;
		16'b1111000001000110 : data_out =  24'b000000000000001000111101;
		16'b1111000001001000 : data_out =  24'b000000000000001000111110;
		16'b1111000001001010 : data_out =  24'b000000000000001000111110;
		16'b1111000001001100 : data_out =  24'b000000000000001000111111;
		16'b1111000001001110 : data_out =  24'b000000000000001000111111;
		16'b1111000001010000 : data_out =  24'b000000000000001001000000;
		16'b1111000001010010 : data_out =  24'b000000000000001001000000;
		16'b1111000001010100 : data_out =  24'b000000000000001001000001;
		16'b1111000001010111 : data_out =  24'b000000000000001001000010;
		16'b1111000001011001 : data_out =  24'b000000000000001001000010;
		16'b1111000001011011 : data_out =  24'b000000000000001001000011;
		16'b1111000001011101 : data_out =  24'b000000000000001001000011;
		16'b1111000001011111 : data_out =  24'b000000000000001001000100;
		16'b1111000001100001 : data_out =  24'b000000000000001001000101;
		16'b1111000001100011 : data_out =  24'b000000000000001001000101;
		16'b1111000001100101 : data_out =  24'b000000000000001001000110;
		16'b1111000001100111 : data_out =  24'b000000000000001001000110;
		16'b1111000001101001 : data_out =  24'b000000000000001001000111;
		16'b1111000001101011 : data_out =  24'b000000000000001001000111;
		16'b1111000001101101 : data_out =  24'b000000000000001001001000;
		16'b1111000001101111 : data_out =  24'b000000000000001001001001;
		16'b1111000001110001 : data_out =  24'b000000000000001001001001;
		16'b1111000001110011 : data_out =  24'b000000000000001001001010;
		16'b1111000001110101 : data_out =  24'b000000000000001001001010;
		16'b1111000001110111 : data_out =  24'b000000000000001001001011;
		16'b1111000001111001 : data_out =  24'b000000000000001001001100;
		16'b1111000001111011 : data_out =  24'b000000000000001001001100;
		16'b1111000001111101 : data_out =  24'b000000000000001001001101;
		16'b1111000001111111 : data_out =  24'b000000000000001001001101;
		16'b1111000010000010 : data_out =  24'b000000000000001001001110;
		16'b1111000010000100 : data_out =  24'b000000000000001001001110;
		16'b1111000010000110 : data_out =  24'b000000000000001001001111;
		16'b1111000010001000 : data_out =  24'b000000000000001001010000;
		16'b1111000010001010 : data_out =  24'b000000000000001001010000;
		16'b1111000010001100 : data_out =  24'b000000000000001001010001;
		16'b1111000010001110 : data_out =  24'b000000000000001001010001;
		16'b1111000010010000 : data_out =  24'b000000000000001001010010;
		16'b1111000010010010 : data_out =  24'b000000000000001001010011;
		16'b1111000010010100 : data_out =  24'b000000000000001001010011;
		16'b1111000010010110 : data_out =  24'b000000000000001001010100;
		16'b1111000010011000 : data_out =  24'b000000000000001001010100;
		16'b1111000010011010 : data_out =  24'b000000000000001001010101;
		16'b1111000010011100 : data_out =  24'b000000000000001001010110;
		16'b1111000010011110 : data_out =  24'b000000000000001001010110;
		16'b1111000010100000 : data_out =  24'b000000000000001001010111;
		16'b1111000010100010 : data_out =  24'b000000000000001001010111;
		16'b1111000010100100 : data_out =  24'b000000000000001001011000;
		16'b1111000010100110 : data_out =  24'b000000000000001001011001;
		16'b1111000010101000 : data_out =  24'b000000000000001001011001;
		16'b1111000010101010 : data_out =  24'b000000000000001001011010;
		16'b1111000010101101 : data_out =  24'b000000000000001001011010;
		16'b1111000010101111 : data_out =  24'b000000000000001001011011;
		16'b1111000010110001 : data_out =  24'b000000000000001001011100;
		16'b1111000010110011 : data_out =  24'b000000000000001001011100;
		16'b1111000010110101 : data_out =  24'b000000000000001001011101;
		16'b1111000010110111 : data_out =  24'b000000000000001001011101;
		16'b1111000010111001 : data_out =  24'b000000000000001001011110;
		16'b1111000010111011 : data_out =  24'b000000000000001001011111;
		16'b1111000010111101 : data_out =  24'b000000000000001001011111;
		16'b1111000010111111 : data_out =  24'b000000000000001001100000;
		16'b1111000011000001 : data_out =  24'b000000000000001001100000;
		16'b1111000011000011 : data_out =  24'b000000000000001001100001;
		16'b1111000011000101 : data_out =  24'b000000000000001001100010;
		16'b1111000011000111 : data_out =  24'b000000000000001001100010;
		16'b1111000011001001 : data_out =  24'b000000000000001001100011;
		16'b1111000011001011 : data_out =  24'b000000000000001001100100;
		16'b1111000011001101 : data_out =  24'b000000000000001001100100;
		16'b1111000011001111 : data_out =  24'b000000000000001001100101;
		16'b1111000011010001 : data_out =  24'b000000000000001001100101;
		16'b1111000011010011 : data_out =  24'b000000000000001001100110;
		16'b1111000011010101 : data_out =  24'b000000000000001001100111;
		16'b1111000011011000 : data_out =  24'b000000000000001001100111;
		16'b1111000011011010 : data_out =  24'b000000000000001001101000;
		16'b1111000011011100 : data_out =  24'b000000000000001001101000;
		16'b1111000011011110 : data_out =  24'b000000000000001001101001;
		16'b1111000011100000 : data_out =  24'b000000000000001001101010;
		16'b1111000011100010 : data_out =  24'b000000000000001001101010;
		16'b1111000011100100 : data_out =  24'b000000000000001001101011;
		16'b1111000011100110 : data_out =  24'b000000000000001001101100;
		16'b1111000011101000 : data_out =  24'b000000000000001001101100;
		16'b1111000011101010 : data_out =  24'b000000000000001001101101;
		16'b1111000011101100 : data_out =  24'b000000000000001001101101;
		16'b1111000011101110 : data_out =  24'b000000000000001001101110;
		16'b1111000011110000 : data_out =  24'b000000000000001001101111;
		16'b1111000011110010 : data_out =  24'b000000000000001001101111;
		16'b1111000011110100 : data_out =  24'b000000000000001001110000;
		16'b1111000011110110 : data_out =  24'b000000000000001001110001;
		16'b1111000011111000 : data_out =  24'b000000000000001001110001;
		16'b1111000011111010 : data_out =  24'b000000000000001001110010;
		16'b1111000011111100 : data_out =  24'b000000000000001001110010;
		16'b1111000011111110 : data_out =  24'b000000000000001001110011;
		16'b1111000100000001 : data_out =  24'b000000000000001001110100;
		16'b1111000100000011 : data_out =  24'b000000000000001001110100;
		16'b1111000100000101 : data_out =  24'b000000000000001001110101;
		16'b1111000100000111 : data_out =  24'b000000000000001001110110;
		16'b1111000100001001 : data_out =  24'b000000000000001001110110;
		16'b1111000100001011 : data_out =  24'b000000000000001001110111;
		16'b1111000100001101 : data_out =  24'b000000000000001001110111;
		16'b1111000100001111 : data_out =  24'b000000000000001001111000;
		16'b1111000100010001 : data_out =  24'b000000000000001001111001;
		16'b1111000100010011 : data_out =  24'b000000000000001001111001;
		16'b1111000100010101 : data_out =  24'b000000000000001001111010;
		16'b1111000100010111 : data_out =  24'b000000000000001001111011;
		16'b1111000100011001 : data_out =  24'b000000000000001001111011;
		16'b1111000100011011 : data_out =  24'b000000000000001001111100;
		16'b1111000100011101 : data_out =  24'b000000000000001001111100;
		16'b1111000100011111 : data_out =  24'b000000000000001001111101;
		16'b1111000100100001 : data_out =  24'b000000000000001001111110;
		16'b1111000100100011 : data_out =  24'b000000000000001001111110;
		16'b1111000100100101 : data_out =  24'b000000000000001001111111;
		16'b1111000100100111 : data_out =  24'b000000000000001010000000;
		16'b1111000100101001 : data_out =  24'b000000000000001010000000;
		16'b1111000100101100 : data_out =  24'b000000000000001010000001;
		16'b1111000100101110 : data_out =  24'b000000000000001010000010;
		16'b1111000100110000 : data_out =  24'b000000000000001010000010;
		16'b1111000100110010 : data_out =  24'b000000000000001010000011;
		16'b1111000100110100 : data_out =  24'b000000000000001010000100;
		16'b1111000100110110 : data_out =  24'b000000000000001010000100;
		16'b1111000100111000 : data_out =  24'b000000000000001010000101;
		16'b1111000100111010 : data_out =  24'b000000000000001010000101;
		16'b1111000100111100 : data_out =  24'b000000000000001010000110;
		16'b1111000100111110 : data_out =  24'b000000000000001010000111;
		16'b1111000101000000 : data_out =  24'b000000000000001010000111;
		16'b1111000101000010 : data_out =  24'b000000000000001010001000;
		16'b1111000101000100 : data_out =  24'b000000000000001010001001;
		16'b1111000101000110 : data_out =  24'b000000000000001010001001;
		16'b1111000101001000 : data_out =  24'b000000000000001010001010;
		16'b1111000101001010 : data_out =  24'b000000000000001010001011;
		16'b1111000101001100 : data_out =  24'b000000000000001010001011;
		16'b1111000101001110 : data_out =  24'b000000000000001010001100;
		16'b1111000101010000 : data_out =  24'b000000000000001010001101;
		16'b1111000101010010 : data_out =  24'b000000000000001010001101;
		16'b1111000101010100 : data_out =  24'b000000000000001010001110;
		16'b1111000101010111 : data_out =  24'b000000000000001010001111;
		16'b1111000101011001 : data_out =  24'b000000000000001010001111;
		16'b1111000101011011 : data_out =  24'b000000000000001010010000;
		16'b1111000101011101 : data_out =  24'b000000000000001010010001;
		16'b1111000101011111 : data_out =  24'b000000000000001010010001;
		16'b1111000101100001 : data_out =  24'b000000000000001010010010;
		16'b1111000101100011 : data_out =  24'b000000000000001010010011;
		16'b1111000101100101 : data_out =  24'b000000000000001010010011;
		16'b1111000101100111 : data_out =  24'b000000000000001010010100;
		16'b1111000101101001 : data_out =  24'b000000000000001010010101;
		16'b1111000101101011 : data_out =  24'b000000000000001010010101;
		16'b1111000101101101 : data_out =  24'b000000000000001010010110;
		16'b1111000101101111 : data_out =  24'b000000000000001010010110;
		16'b1111000101110001 : data_out =  24'b000000000000001010010111;
		16'b1111000101110011 : data_out =  24'b000000000000001010011000;
		16'b1111000101110101 : data_out =  24'b000000000000001010011000;
		16'b1111000101110111 : data_out =  24'b000000000000001010011001;
		16'b1111000101111001 : data_out =  24'b000000000000001010011010;
		16'b1111000101111011 : data_out =  24'b000000000000001010011010;
		16'b1111000101111101 : data_out =  24'b000000000000001010011011;
		16'b1111000101111111 : data_out =  24'b000000000000001010011100;
		16'b1111000110000010 : data_out =  24'b000000000000001010011100;
		16'b1111000110000100 : data_out =  24'b000000000000001010011101;
		16'b1111000110000110 : data_out =  24'b000000000000001010011110;
		16'b1111000110001000 : data_out =  24'b000000000000001010011110;
		16'b1111000110001010 : data_out =  24'b000000000000001010011111;
		16'b1111000110001100 : data_out =  24'b000000000000001010100000;
		16'b1111000110001110 : data_out =  24'b000000000000001010100001;
		16'b1111000110010000 : data_out =  24'b000000000000001010100001;
		16'b1111000110010010 : data_out =  24'b000000000000001010100010;
		16'b1111000110010100 : data_out =  24'b000000000000001010100011;
		16'b1111000110010110 : data_out =  24'b000000000000001010100011;
		16'b1111000110011000 : data_out =  24'b000000000000001010100100;
		16'b1111000110011010 : data_out =  24'b000000000000001010100101;
		16'b1111000110011100 : data_out =  24'b000000000000001010100101;
		16'b1111000110011110 : data_out =  24'b000000000000001010100110;
		16'b1111000110100000 : data_out =  24'b000000000000001010100111;
		16'b1111000110100010 : data_out =  24'b000000000000001010100111;
		16'b1111000110100100 : data_out =  24'b000000000000001010101000;
		16'b1111000110100110 : data_out =  24'b000000000000001010101001;
		16'b1111000110101000 : data_out =  24'b000000000000001010101001;
		16'b1111000110101010 : data_out =  24'b000000000000001010101010;
		16'b1111000110101101 : data_out =  24'b000000000000001010101011;
		16'b1111000110101111 : data_out =  24'b000000000000001010101011;
		16'b1111000110110001 : data_out =  24'b000000000000001010101100;
		16'b1111000110110011 : data_out =  24'b000000000000001010101101;
		16'b1111000110110101 : data_out =  24'b000000000000001010101101;
		16'b1111000110110111 : data_out =  24'b000000000000001010101110;
		16'b1111000110111001 : data_out =  24'b000000000000001010101111;
		16'b1111000110111011 : data_out =  24'b000000000000001010101111;
		16'b1111000110111101 : data_out =  24'b000000000000001010110000;
		16'b1111000110111111 : data_out =  24'b000000000000001010110001;
		16'b1111000111000001 : data_out =  24'b000000000000001010110010;
		16'b1111000111000011 : data_out =  24'b000000000000001010110010;
		16'b1111000111000101 : data_out =  24'b000000000000001010110011;
		16'b1111000111000111 : data_out =  24'b000000000000001010110100;
		16'b1111000111001001 : data_out =  24'b000000000000001010110100;
		16'b1111000111001011 : data_out =  24'b000000000000001010110101;
		16'b1111000111001101 : data_out =  24'b000000000000001010110110;
		16'b1111000111001111 : data_out =  24'b000000000000001010110110;
		16'b1111000111010001 : data_out =  24'b000000000000001010110111;
		16'b1111000111010011 : data_out =  24'b000000000000001010111000;
		16'b1111000111010101 : data_out =  24'b000000000000001010111000;
		16'b1111000111011000 : data_out =  24'b000000000000001010111001;
		16'b1111000111011010 : data_out =  24'b000000000000001010111010;
		16'b1111000111011100 : data_out =  24'b000000000000001010111011;
		16'b1111000111011110 : data_out =  24'b000000000000001010111011;
		16'b1111000111100000 : data_out =  24'b000000000000001010111100;
		16'b1111000111100010 : data_out =  24'b000000000000001010111101;
		16'b1111000111100100 : data_out =  24'b000000000000001010111101;
		16'b1111000111100110 : data_out =  24'b000000000000001010111110;
		16'b1111000111101000 : data_out =  24'b000000000000001010111111;
		16'b1111000111101010 : data_out =  24'b000000000000001010111111;
		16'b1111000111101100 : data_out =  24'b000000000000001011000000;
		16'b1111000111101110 : data_out =  24'b000000000000001011000001;
		16'b1111000111110000 : data_out =  24'b000000000000001011000010;
		16'b1111000111110010 : data_out =  24'b000000000000001011000010;
		16'b1111000111110100 : data_out =  24'b000000000000001011000011;
		16'b1111000111110110 : data_out =  24'b000000000000001011000100;
		16'b1111000111111000 : data_out =  24'b000000000000001011000100;
		16'b1111000111111010 : data_out =  24'b000000000000001011000101;
		16'b1111000111111100 : data_out =  24'b000000000000001011000110;
		16'b1111000111111110 : data_out =  24'b000000000000001011000111;
		16'b1111001000000001 : data_out =  24'b000000000000001011000111;
		16'b1111001000000011 : data_out =  24'b000000000000001011001000;
		16'b1111001000000101 : data_out =  24'b000000000000001011001001;
		16'b1111001000000111 : data_out =  24'b000000000000001011001001;
		16'b1111001000001001 : data_out =  24'b000000000000001011001010;
		16'b1111001000001011 : data_out =  24'b000000000000001011001011;
		16'b1111001000001101 : data_out =  24'b000000000000001011001100;
		16'b1111001000001111 : data_out =  24'b000000000000001011001100;
		16'b1111001000010001 : data_out =  24'b000000000000001011001101;
		16'b1111001000010011 : data_out =  24'b000000000000001011001110;
		16'b1111001000010101 : data_out =  24'b000000000000001011001110;
		16'b1111001000010111 : data_out =  24'b000000000000001011001111;
		16'b1111001000011001 : data_out =  24'b000000000000001011010000;
		16'b1111001000011011 : data_out =  24'b000000000000001011010001;
		16'b1111001000011101 : data_out =  24'b000000000000001011010001;
		16'b1111001000011111 : data_out =  24'b000000000000001011010010;
		16'b1111001000100001 : data_out =  24'b000000000000001011010011;
		16'b1111001000100011 : data_out =  24'b000000000000001011010011;
		16'b1111001000100101 : data_out =  24'b000000000000001011010100;
		16'b1111001000100111 : data_out =  24'b000000000000001011010101;
		16'b1111001000101001 : data_out =  24'b000000000000001011010110;
		16'b1111001000101100 : data_out =  24'b000000000000001011010110;
		16'b1111001000101110 : data_out =  24'b000000000000001011010111;
		16'b1111001000110000 : data_out =  24'b000000000000001011011000;
		16'b1111001000110010 : data_out =  24'b000000000000001011011001;
		16'b1111001000110100 : data_out =  24'b000000000000001011011001;
		16'b1111001000110110 : data_out =  24'b000000000000001011011010;
		16'b1111001000111000 : data_out =  24'b000000000000001011011011;
		16'b1111001000111010 : data_out =  24'b000000000000001011011011;
		16'b1111001000111100 : data_out =  24'b000000000000001011011100;
		16'b1111001000111110 : data_out =  24'b000000000000001011011101;
		16'b1111001001000000 : data_out =  24'b000000000000001011011110;
		16'b1111001001000010 : data_out =  24'b000000000000001011011110;
		16'b1111001001000100 : data_out =  24'b000000000000001011011111;
		16'b1111001001000110 : data_out =  24'b000000000000001011100000;
		16'b1111001001001000 : data_out =  24'b000000000000001011100001;
		16'b1111001001001010 : data_out =  24'b000000000000001011100001;
		16'b1111001001001100 : data_out =  24'b000000000000001011100010;
		16'b1111001001001110 : data_out =  24'b000000000000001011100011;
		16'b1111001001010000 : data_out =  24'b000000000000001011100100;
		16'b1111001001010010 : data_out =  24'b000000000000001011100100;
		16'b1111001001010100 : data_out =  24'b000000000000001011100101;
		16'b1111001001010111 : data_out =  24'b000000000000001011100110;
		16'b1111001001011001 : data_out =  24'b000000000000001011100111;
		16'b1111001001011011 : data_out =  24'b000000000000001011100111;
		16'b1111001001011101 : data_out =  24'b000000000000001011101000;
		16'b1111001001011111 : data_out =  24'b000000000000001011101001;
		16'b1111001001100001 : data_out =  24'b000000000000001011101010;
		16'b1111001001100011 : data_out =  24'b000000000000001011101010;
		16'b1111001001100101 : data_out =  24'b000000000000001011101011;
		16'b1111001001100111 : data_out =  24'b000000000000001011101100;
		16'b1111001001101001 : data_out =  24'b000000000000001011101101;
		16'b1111001001101011 : data_out =  24'b000000000000001011101101;
		16'b1111001001101101 : data_out =  24'b000000000000001011101110;
		16'b1111001001101111 : data_out =  24'b000000000000001011101111;
		16'b1111001001110001 : data_out =  24'b000000000000001011110000;
		16'b1111001001110011 : data_out =  24'b000000000000001011110000;
		16'b1111001001110101 : data_out =  24'b000000000000001011110001;
		16'b1111001001110111 : data_out =  24'b000000000000001011110010;
		16'b1111001001111001 : data_out =  24'b000000000000001011110011;
		16'b1111001001111011 : data_out =  24'b000000000000001011110011;
		16'b1111001001111101 : data_out =  24'b000000000000001011110100;
		16'b1111001001111111 : data_out =  24'b000000000000001011110101;
		16'b1111001010000010 : data_out =  24'b000000000000001011110110;
		16'b1111001010000100 : data_out =  24'b000000000000001011110110;
		16'b1111001010000110 : data_out =  24'b000000000000001011110111;
		16'b1111001010001000 : data_out =  24'b000000000000001011111000;
		16'b1111001010001010 : data_out =  24'b000000000000001011111001;
		16'b1111001010001100 : data_out =  24'b000000000000001011111001;
		16'b1111001010001110 : data_out =  24'b000000000000001011111010;
		16'b1111001010010000 : data_out =  24'b000000000000001011111011;
		16'b1111001010010010 : data_out =  24'b000000000000001011111100;
		16'b1111001010010100 : data_out =  24'b000000000000001011111100;
		16'b1111001010010110 : data_out =  24'b000000000000001011111101;
		16'b1111001010011000 : data_out =  24'b000000000000001011111110;
		16'b1111001010011010 : data_out =  24'b000000000000001011111111;
		16'b1111001010011100 : data_out =  24'b000000000000001011111111;
		16'b1111001010011110 : data_out =  24'b000000000000001100000000;
		16'b1111001010100000 : data_out =  24'b000000000000001100000001;
		16'b1111001010100010 : data_out =  24'b000000000000001100000010;
		16'b1111001010100100 : data_out =  24'b000000000000001100000011;
		16'b1111001010100110 : data_out =  24'b000000000000001100000011;
		16'b1111001010101000 : data_out =  24'b000000000000001100000100;
		16'b1111001010101010 : data_out =  24'b000000000000001100000101;
		16'b1111001010101101 : data_out =  24'b000000000000001100000110;
		16'b1111001010101111 : data_out =  24'b000000000000001100000110;
		16'b1111001010110001 : data_out =  24'b000000000000001100000111;
		16'b1111001010110011 : data_out =  24'b000000000000001100001000;
		16'b1111001010110101 : data_out =  24'b000000000000001100001001;
		16'b1111001010110111 : data_out =  24'b000000000000001100001010;
		16'b1111001010111001 : data_out =  24'b000000000000001100001010;
		16'b1111001010111011 : data_out =  24'b000000000000001100001011;
		16'b1111001010111101 : data_out =  24'b000000000000001100001100;
		16'b1111001010111111 : data_out =  24'b000000000000001100001101;
		16'b1111001011000001 : data_out =  24'b000000000000001100001101;
		16'b1111001011000011 : data_out =  24'b000000000000001100001110;
		16'b1111001011000101 : data_out =  24'b000000000000001100001111;
		16'b1111001011000111 : data_out =  24'b000000000000001100010000;
		16'b1111001011001001 : data_out =  24'b000000000000001100010001;
		16'b1111001011001011 : data_out =  24'b000000000000001100010001;
		16'b1111001011001101 : data_out =  24'b000000000000001100010010;
		16'b1111001011001111 : data_out =  24'b000000000000001100010011;
		16'b1111001011010001 : data_out =  24'b000000000000001100010100;
		16'b1111001011010011 : data_out =  24'b000000000000001100010100;
		16'b1111001011010101 : data_out =  24'b000000000000001100010101;
		16'b1111001011011000 : data_out =  24'b000000000000001100010110;
		16'b1111001011011010 : data_out =  24'b000000000000001100010111;
		16'b1111001011011100 : data_out =  24'b000000000000001100011000;
		16'b1111001011011110 : data_out =  24'b000000000000001100011000;
		16'b1111001011100000 : data_out =  24'b000000000000001100011001;
		16'b1111001011100010 : data_out =  24'b000000000000001100011010;
		16'b1111001011100100 : data_out =  24'b000000000000001100011011;
		16'b1111001011100110 : data_out =  24'b000000000000001100011100;
		16'b1111001011101000 : data_out =  24'b000000000000001100011100;
		16'b1111001011101010 : data_out =  24'b000000000000001100011101;
		16'b1111001011101100 : data_out =  24'b000000000000001100011110;
		16'b1111001011101110 : data_out =  24'b000000000000001100011111;
		16'b1111001011110000 : data_out =  24'b000000000000001100100000;
		16'b1111001011110010 : data_out =  24'b000000000000001100100000;
		16'b1111001011110100 : data_out =  24'b000000000000001100100001;
		16'b1111001011110110 : data_out =  24'b000000000000001100100010;
		16'b1111001011111000 : data_out =  24'b000000000000001100100011;
		16'b1111001011111010 : data_out =  24'b000000000000001100100100;
		16'b1111001011111100 : data_out =  24'b000000000000001100100100;
		16'b1111001011111110 : data_out =  24'b000000000000001100100101;
		16'b1111001100000001 : data_out =  24'b000000000000001100100110;
		16'b1111001100000011 : data_out =  24'b000000000000001100100111;
		16'b1111001100000101 : data_out =  24'b000000000000001100101000;
		16'b1111001100000111 : data_out =  24'b000000000000001100101000;
		16'b1111001100001001 : data_out =  24'b000000000000001100101001;
		16'b1111001100001011 : data_out =  24'b000000000000001100101010;
		16'b1111001100001101 : data_out =  24'b000000000000001100101011;
		16'b1111001100001111 : data_out =  24'b000000000000001100101100;
		16'b1111001100010001 : data_out =  24'b000000000000001100101101;
		16'b1111001100010011 : data_out =  24'b000000000000001100101101;
		16'b1111001100010101 : data_out =  24'b000000000000001100101110;
		16'b1111001100010111 : data_out =  24'b000000000000001100101111;
		16'b1111001100011001 : data_out =  24'b000000000000001100110000;
		16'b1111001100011011 : data_out =  24'b000000000000001100110001;
		16'b1111001100011101 : data_out =  24'b000000000000001100110001;
		16'b1111001100011111 : data_out =  24'b000000000000001100110010;
		16'b1111001100100001 : data_out =  24'b000000000000001100110011;
		16'b1111001100100011 : data_out =  24'b000000000000001100110100;
		16'b1111001100100101 : data_out =  24'b000000000000001100110101;
		16'b1111001100100111 : data_out =  24'b000000000000001100110110;
		16'b1111001100101001 : data_out =  24'b000000000000001100110110;
		16'b1111001100101100 : data_out =  24'b000000000000001100110111;
		16'b1111001100101110 : data_out =  24'b000000000000001100111000;
		16'b1111001100110000 : data_out =  24'b000000000000001100111001;
		16'b1111001100110010 : data_out =  24'b000000000000001100111010;
		16'b1111001100110100 : data_out =  24'b000000000000001100111010;
		16'b1111001100110110 : data_out =  24'b000000000000001100111011;
		16'b1111001100111000 : data_out =  24'b000000000000001100111100;
		16'b1111001100111010 : data_out =  24'b000000000000001100111101;
		16'b1111001100111100 : data_out =  24'b000000000000001100111110;
		16'b1111001100111110 : data_out =  24'b000000000000001100111111;
		16'b1111001101000000 : data_out =  24'b000000000000001100111111;
		16'b1111001101000010 : data_out =  24'b000000000000001101000000;
		16'b1111001101000100 : data_out =  24'b000000000000001101000001;
		16'b1111001101000110 : data_out =  24'b000000000000001101000010;
		16'b1111001101001000 : data_out =  24'b000000000000001101000011;
		16'b1111001101001010 : data_out =  24'b000000000000001101000100;
		16'b1111001101001100 : data_out =  24'b000000000000001101000100;
		16'b1111001101001110 : data_out =  24'b000000000000001101000101;
		16'b1111001101010000 : data_out =  24'b000000000000001101000110;
		16'b1111001101010010 : data_out =  24'b000000000000001101000111;
		16'b1111001101010100 : data_out =  24'b000000000000001101001000;
		16'b1111001101010111 : data_out =  24'b000000000000001101001001;
		16'b1111001101011001 : data_out =  24'b000000000000001101001001;
		16'b1111001101011011 : data_out =  24'b000000000000001101001010;
		16'b1111001101011101 : data_out =  24'b000000000000001101001011;
		16'b1111001101011111 : data_out =  24'b000000000000001101001100;
		16'b1111001101100001 : data_out =  24'b000000000000001101001101;
		16'b1111001101100011 : data_out =  24'b000000000000001101001110;
		16'b1111001101100101 : data_out =  24'b000000000000001101001111;
		16'b1111001101100111 : data_out =  24'b000000000000001101001111;
		16'b1111001101101001 : data_out =  24'b000000000000001101010000;
		16'b1111001101101011 : data_out =  24'b000000000000001101010001;
		16'b1111001101101101 : data_out =  24'b000000000000001101010010;
		16'b1111001101101111 : data_out =  24'b000000000000001101010011;
		16'b1111001101110001 : data_out =  24'b000000000000001101010100;
		16'b1111001101110011 : data_out =  24'b000000000000001101010101;
		16'b1111001101110101 : data_out =  24'b000000000000001101010101;
		16'b1111001101110111 : data_out =  24'b000000000000001101010110;
		16'b1111001101111001 : data_out =  24'b000000000000001101010111;
		16'b1111001101111011 : data_out =  24'b000000000000001101011000;
		16'b1111001101111101 : data_out =  24'b000000000000001101011001;
		16'b1111001101111111 : data_out =  24'b000000000000001101011010;
		16'b1111001110000010 : data_out =  24'b000000000000001101011010;
		16'b1111001110000100 : data_out =  24'b000000000000001101011011;
		16'b1111001110000110 : data_out =  24'b000000000000001101011100;
		16'b1111001110001000 : data_out =  24'b000000000000001101011101;
		16'b1111001110001010 : data_out =  24'b000000000000001101011110;
		16'b1111001110001100 : data_out =  24'b000000000000001101011111;
		16'b1111001110001110 : data_out =  24'b000000000000001101100000;
		16'b1111001110010000 : data_out =  24'b000000000000001101100001;
		16'b1111001110010010 : data_out =  24'b000000000000001101100001;
		16'b1111001110010100 : data_out =  24'b000000000000001101100010;
		16'b1111001110010110 : data_out =  24'b000000000000001101100011;
		16'b1111001110011000 : data_out =  24'b000000000000001101100100;
		16'b1111001110011010 : data_out =  24'b000000000000001101100101;
		16'b1111001110011100 : data_out =  24'b000000000000001101100110;
		16'b1111001110011110 : data_out =  24'b000000000000001101100111;
		16'b1111001110100000 : data_out =  24'b000000000000001101100111;
		16'b1111001110100010 : data_out =  24'b000000000000001101101000;
		16'b1111001110100100 : data_out =  24'b000000000000001101101001;
		16'b1111001110100110 : data_out =  24'b000000000000001101101010;
		16'b1111001110101000 : data_out =  24'b000000000000001101101011;
		16'b1111001110101010 : data_out =  24'b000000000000001101101100;
		16'b1111001110101101 : data_out =  24'b000000000000001101101101;
		16'b1111001110101111 : data_out =  24'b000000000000001101101110;
		16'b1111001110110001 : data_out =  24'b000000000000001101101110;
		16'b1111001110110011 : data_out =  24'b000000000000001101101111;
		16'b1111001110110101 : data_out =  24'b000000000000001101110000;
		16'b1111001110110111 : data_out =  24'b000000000000001101110001;
		16'b1111001110111001 : data_out =  24'b000000000000001101110010;
		16'b1111001110111011 : data_out =  24'b000000000000001101110011;
		16'b1111001110111101 : data_out =  24'b000000000000001101110100;
		16'b1111001110111111 : data_out =  24'b000000000000001101110101;
		16'b1111001111000001 : data_out =  24'b000000000000001101110110;
		16'b1111001111000011 : data_out =  24'b000000000000001101110110;
		16'b1111001111000101 : data_out =  24'b000000000000001101110111;
		16'b1111001111000111 : data_out =  24'b000000000000001101111000;
		16'b1111001111001001 : data_out =  24'b000000000000001101111001;
		16'b1111001111001011 : data_out =  24'b000000000000001101111010;
		16'b1111001111001101 : data_out =  24'b000000000000001101111011;
		16'b1111001111001111 : data_out =  24'b000000000000001101111100;
		16'b1111001111010001 : data_out =  24'b000000000000001101111101;
		16'b1111001111010011 : data_out =  24'b000000000000001101111110;
		16'b1111001111010101 : data_out =  24'b000000000000001101111110;
		16'b1111001111011000 : data_out =  24'b000000000000001101111111;
		16'b1111001111011010 : data_out =  24'b000000000000001110000000;
		16'b1111001111011100 : data_out =  24'b000000000000001110000001;
		16'b1111001111011110 : data_out =  24'b000000000000001110000010;
		16'b1111001111100000 : data_out =  24'b000000000000001110000011;
		16'b1111001111100010 : data_out =  24'b000000000000001110000100;
		16'b1111001111100100 : data_out =  24'b000000000000001110000101;
		16'b1111001111100110 : data_out =  24'b000000000000001110000110;
		16'b1111001111101000 : data_out =  24'b000000000000001110000111;
		16'b1111001111101010 : data_out =  24'b000000000000001110000111;
		16'b1111001111101100 : data_out =  24'b000000000000001110001000;
		16'b1111001111101110 : data_out =  24'b000000000000001110001001;
		16'b1111001111110000 : data_out =  24'b000000000000001110001010;
		16'b1111001111110010 : data_out =  24'b000000000000001110001011;
		16'b1111001111110100 : data_out =  24'b000000000000001110001100;
		16'b1111001111110110 : data_out =  24'b000000000000001110001101;
		16'b1111001111111000 : data_out =  24'b000000000000001110001110;
		16'b1111001111111010 : data_out =  24'b000000000000001110001111;
		16'b1111001111111100 : data_out =  24'b000000000000001110010000;
		16'b1111001111111110 : data_out =  24'b000000000000001110010001;
		16'b1111010000000001 : data_out =  24'b000000000000001110010001;
		16'b1111010000000011 : data_out =  24'b000000000000001110010010;
		16'b1111010000000101 : data_out =  24'b000000000000001110010011;
		16'b1111010000000111 : data_out =  24'b000000000000001110010100;
		16'b1111010000001001 : data_out =  24'b000000000000001110010101;
		16'b1111010000001011 : data_out =  24'b000000000000001110010110;
		16'b1111010000001101 : data_out =  24'b000000000000001110010111;
		16'b1111010000001111 : data_out =  24'b000000000000001110011000;
		16'b1111010000010001 : data_out =  24'b000000000000001110011001;
		16'b1111010000010011 : data_out =  24'b000000000000001110011010;
		16'b1111010000010101 : data_out =  24'b000000000000001110011011;
		16'b1111010000010111 : data_out =  24'b000000000000001110011100;
		16'b1111010000011001 : data_out =  24'b000000000000001110011100;
		16'b1111010000011011 : data_out =  24'b000000000000001110011101;
		16'b1111010000011101 : data_out =  24'b000000000000001110011110;
		16'b1111010000011111 : data_out =  24'b000000000000001110011111;
		16'b1111010000100001 : data_out =  24'b000000000000001110100000;
		16'b1111010000100011 : data_out =  24'b000000000000001110100001;
		16'b1111010000100101 : data_out =  24'b000000000000001110100010;
		16'b1111010000100111 : data_out =  24'b000000000000001110100011;
		16'b1111010000101001 : data_out =  24'b000000000000001110100100;
		16'b1111010000101100 : data_out =  24'b000000000000001110100101;
		16'b1111010000101110 : data_out =  24'b000000000000001110100110;
		16'b1111010000110000 : data_out =  24'b000000000000001110100111;
		16'b1111010000110010 : data_out =  24'b000000000000001110101000;
		16'b1111010000110100 : data_out =  24'b000000000000001110101001;
		16'b1111010000110110 : data_out =  24'b000000000000001110101010;
		16'b1111010000111000 : data_out =  24'b000000000000001110101010;
		16'b1111010000111010 : data_out =  24'b000000000000001110101011;
		16'b1111010000111100 : data_out =  24'b000000000000001110101100;
		16'b1111010000111110 : data_out =  24'b000000000000001110101101;
		16'b1111010001000000 : data_out =  24'b000000000000001110101110;
		16'b1111010001000010 : data_out =  24'b000000000000001110101111;
		16'b1111010001000100 : data_out =  24'b000000000000001110110000;
		16'b1111010001000110 : data_out =  24'b000000000000001110110001;
		16'b1111010001001000 : data_out =  24'b000000000000001110110010;
		16'b1111010001001010 : data_out =  24'b000000000000001110110011;
		16'b1111010001001100 : data_out =  24'b000000000000001110110100;
		16'b1111010001001110 : data_out =  24'b000000000000001110110101;
		16'b1111010001010000 : data_out =  24'b000000000000001110110110;
		16'b1111010001010010 : data_out =  24'b000000000000001110110111;
		16'b1111010001010100 : data_out =  24'b000000000000001110111000;
		16'b1111010001010111 : data_out =  24'b000000000000001110111001;
		16'b1111010001011001 : data_out =  24'b000000000000001110111010;
		16'b1111010001011011 : data_out =  24'b000000000000001110111011;
		16'b1111010001011101 : data_out =  24'b000000000000001110111100;
		16'b1111010001011111 : data_out =  24'b000000000000001110111100;
		16'b1111010001100001 : data_out =  24'b000000000000001110111101;
		16'b1111010001100011 : data_out =  24'b000000000000001110111110;
		16'b1111010001100101 : data_out =  24'b000000000000001110111111;
		16'b1111010001100111 : data_out =  24'b000000000000001111000000;
		16'b1111010001101001 : data_out =  24'b000000000000001111000001;
		16'b1111010001101011 : data_out =  24'b000000000000001111000010;
		16'b1111010001101101 : data_out =  24'b000000000000001111000011;
		16'b1111010001101111 : data_out =  24'b000000000000001111000100;
		16'b1111010001110001 : data_out =  24'b000000000000001111000101;
		16'b1111010001110011 : data_out =  24'b000000000000001111000110;
		16'b1111010001110101 : data_out =  24'b000000000000001111000111;
		16'b1111010001110111 : data_out =  24'b000000000000001111001000;
		16'b1111010001111001 : data_out =  24'b000000000000001111001001;
		16'b1111010001111011 : data_out =  24'b000000000000001111001010;
		16'b1111010001111101 : data_out =  24'b000000000000001111001011;
		16'b1111010001111111 : data_out =  24'b000000000000001111001100;
		16'b1111010010000010 : data_out =  24'b000000000000001111001101;
		16'b1111010010000100 : data_out =  24'b000000000000001111001110;
		16'b1111010010000110 : data_out =  24'b000000000000001111001111;
		16'b1111010010001000 : data_out =  24'b000000000000001111010000;
		16'b1111010010001010 : data_out =  24'b000000000000001111010001;
		16'b1111010010001100 : data_out =  24'b000000000000001111010010;
		16'b1111010010001110 : data_out =  24'b000000000000001111010011;
		16'b1111010010010000 : data_out =  24'b000000000000001111010100;
		16'b1111010010010010 : data_out =  24'b000000000000001111010101;
		16'b1111010010010100 : data_out =  24'b000000000000001111010110;
		16'b1111010010010110 : data_out =  24'b000000000000001111010111;
		16'b1111010010011000 : data_out =  24'b000000000000001111011000;
		16'b1111010010011010 : data_out =  24'b000000000000001111011001;
		16'b1111010010011100 : data_out =  24'b000000000000001111011010;
		16'b1111010010011110 : data_out =  24'b000000000000001111011011;
		16'b1111010010100000 : data_out =  24'b000000000000001111011100;
		16'b1111010010100010 : data_out =  24'b000000000000001111011101;
		16'b1111010010100100 : data_out =  24'b000000000000001111011110;
		16'b1111010010100110 : data_out =  24'b000000000000001111011111;
		16'b1111010010101000 : data_out =  24'b000000000000001111100000;
		16'b1111010010101010 : data_out =  24'b000000000000001111100001;
		16'b1111010010101101 : data_out =  24'b000000000000001111100010;
		16'b1111010010101111 : data_out =  24'b000000000000001111100011;
		16'b1111010010110001 : data_out =  24'b000000000000001111100100;
		16'b1111010010110011 : data_out =  24'b000000000000001111100101;
		16'b1111010010110101 : data_out =  24'b000000000000001111100110;
		16'b1111010010110111 : data_out =  24'b000000000000001111100111;
		16'b1111010010111001 : data_out =  24'b000000000000001111101000;
		16'b1111010010111011 : data_out =  24'b000000000000001111101001;
		16'b1111010010111101 : data_out =  24'b000000000000001111101010;
		16'b1111010010111111 : data_out =  24'b000000000000001111101011;
		16'b1111010011000001 : data_out =  24'b000000000000001111101100;
		16'b1111010011000011 : data_out =  24'b000000000000001111101101;
		16'b1111010011000101 : data_out =  24'b000000000000001111101110;
		16'b1111010011000111 : data_out =  24'b000000000000001111101111;
		16'b1111010011001001 : data_out =  24'b000000000000001111110000;
		16'b1111010011001011 : data_out =  24'b000000000000001111110001;
		16'b1111010011001101 : data_out =  24'b000000000000001111110010;
		16'b1111010011001111 : data_out =  24'b000000000000001111110011;
		16'b1111010011010001 : data_out =  24'b000000000000001111110100;
		16'b1111010011010011 : data_out =  24'b000000000000001111110101;
		16'b1111010011010101 : data_out =  24'b000000000000001111110110;
		16'b1111010011011000 : data_out =  24'b000000000000001111110111;
		16'b1111010011011010 : data_out =  24'b000000000000001111111000;
		16'b1111010011011100 : data_out =  24'b000000000000001111111001;
		16'b1111010011011110 : data_out =  24'b000000000000001111111010;
		16'b1111010011100000 : data_out =  24'b000000000000001111111011;
		16'b1111010011100010 : data_out =  24'b000000000000001111111100;
		16'b1111010011100100 : data_out =  24'b000000000000001111111101;
		16'b1111010011100110 : data_out =  24'b000000000000001111111110;
		16'b1111010011101000 : data_out =  24'b000000000000001111111111;
		16'b1111010011101010 : data_out =  24'b000000000000010000000000;
		16'b1111010011101100 : data_out =  24'b000000000000010000000001;
		16'b1111010011101110 : data_out =  24'b000000000000010000000010;
		16'b1111010011110000 : data_out =  24'b000000000000010000000011;
		16'b1111010011110010 : data_out =  24'b000000000000010000000100;
		16'b1111010011110100 : data_out =  24'b000000000000010000000101;
		16'b1111010011110110 : data_out =  24'b000000000000010000000110;
		16'b1111010011111000 : data_out =  24'b000000000000010000000111;
		16'b1111010011111010 : data_out =  24'b000000000000010000001000;
		16'b1111010011111100 : data_out =  24'b000000000000010000001001;
		16'b1111010011111110 : data_out =  24'b000000000000010000001010;
		16'b1111010100000001 : data_out =  24'b000000000000010000001011;
		16'b1111010100000011 : data_out =  24'b000000000000010000001100;
		16'b1111010100000101 : data_out =  24'b000000000000010000001101;
		16'b1111010100000111 : data_out =  24'b000000000000010000001110;
		16'b1111010100001001 : data_out =  24'b000000000000010000001111;
		16'b1111010100001011 : data_out =  24'b000000000000010000010000;
		16'b1111010100001101 : data_out =  24'b000000000000010000010001;
		16'b1111010100001111 : data_out =  24'b000000000000010000010010;
		16'b1111010100010001 : data_out =  24'b000000000000010000010011;
		16'b1111010100010011 : data_out =  24'b000000000000010000010100;
		16'b1111010100010101 : data_out =  24'b000000000000010000010110;
		16'b1111010100010111 : data_out =  24'b000000000000010000010111;
		16'b1111010100011001 : data_out =  24'b000000000000010000011000;
		16'b1111010100011011 : data_out =  24'b000000000000010000011001;
		16'b1111010100011101 : data_out =  24'b000000000000010000011010;
		16'b1111010100011111 : data_out =  24'b000000000000010000011011;
		16'b1111010100100001 : data_out =  24'b000000000000010000011100;
		16'b1111010100100011 : data_out =  24'b000000000000010000011101;
		16'b1111010100100101 : data_out =  24'b000000000000010000011110;
		16'b1111010100100111 : data_out =  24'b000000000000010000011111;
		16'b1111010100101001 : data_out =  24'b000000000000010000100000;
		16'b1111010100101100 : data_out =  24'b000000000000010000100001;
		16'b1111010100101110 : data_out =  24'b000000000000010000100010;
		16'b1111010100110000 : data_out =  24'b000000000000010000100011;
		16'b1111010100110010 : data_out =  24'b000000000000010000100100;
		16'b1111010100110100 : data_out =  24'b000000000000010000100101;
		16'b1111010100110110 : data_out =  24'b000000000000010000100110;
		16'b1111010100111000 : data_out =  24'b000000000000010000100111;
		16'b1111010100111010 : data_out =  24'b000000000000010000101001;
		16'b1111010100111100 : data_out =  24'b000000000000010000101010;
		16'b1111010100111110 : data_out =  24'b000000000000010000101011;
		16'b1111010101000000 : data_out =  24'b000000000000010000101100;
		16'b1111010101000010 : data_out =  24'b000000000000010000101101;
		16'b1111010101000100 : data_out =  24'b000000000000010000101110;
		16'b1111010101000110 : data_out =  24'b000000000000010000101111;
		16'b1111010101001000 : data_out =  24'b000000000000010000110000;
		16'b1111010101001010 : data_out =  24'b000000000000010000110001;
		16'b1111010101001100 : data_out =  24'b000000000000010000110010;
		16'b1111010101001110 : data_out =  24'b000000000000010000110011;
		16'b1111010101010000 : data_out =  24'b000000000000010000110100;
		16'b1111010101010010 : data_out =  24'b000000000000010000110101;
		16'b1111010101010100 : data_out =  24'b000000000000010000110110;
		16'b1111010101010111 : data_out =  24'b000000000000010000111000;
		16'b1111010101011001 : data_out =  24'b000000000000010000111001;
		16'b1111010101011011 : data_out =  24'b000000000000010000111010;
		16'b1111010101011101 : data_out =  24'b000000000000010000111011;
		16'b1111010101011111 : data_out =  24'b000000000000010000111100;
		16'b1111010101100001 : data_out =  24'b000000000000010000111101;
		16'b1111010101100011 : data_out =  24'b000000000000010000111110;
		16'b1111010101100101 : data_out =  24'b000000000000010000111111;
		16'b1111010101100111 : data_out =  24'b000000000000010001000000;
		16'b1111010101101001 : data_out =  24'b000000000000010001000001;
		16'b1111010101101011 : data_out =  24'b000000000000010001000010;
		16'b1111010101101101 : data_out =  24'b000000000000010001000100;
		16'b1111010101101111 : data_out =  24'b000000000000010001000101;
		16'b1111010101110001 : data_out =  24'b000000000000010001000110;
		16'b1111010101110011 : data_out =  24'b000000000000010001000111;
		16'b1111010101110101 : data_out =  24'b000000000000010001001000;
		16'b1111010101110111 : data_out =  24'b000000000000010001001001;
		16'b1111010101111001 : data_out =  24'b000000000000010001001010;
		16'b1111010101111011 : data_out =  24'b000000000000010001001011;
		16'b1111010101111101 : data_out =  24'b000000000000010001001100;
		16'b1111010101111111 : data_out =  24'b000000000000010001001101;
		16'b1111010110000010 : data_out =  24'b000000000000010001001110;
		16'b1111010110000100 : data_out =  24'b000000000000010001010000;
		16'b1111010110000110 : data_out =  24'b000000000000010001010001;
		16'b1111010110001000 : data_out =  24'b000000000000010001010010;
		16'b1111010110001010 : data_out =  24'b000000000000010001010011;
		16'b1111010110001100 : data_out =  24'b000000000000010001010100;
		16'b1111010110001110 : data_out =  24'b000000000000010001010101;
		16'b1111010110010000 : data_out =  24'b000000000000010001010110;
		16'b1111010110010010 : data_out =  24'b000000000000010001010111;
		16'b1111010110010100 : data_out =  24'b000000000000010001011000;
		16'b1111010110010110 : data_out =  24'b000000000000010001011010;
		16'b1111010110011000 : data_out =  24'b000000000000010001011011;
		16'b1111010110011010 : data_out =  24'b000000000000010001011100;
		16'b1111010110011100 : data_out =  24'b000000000000010001011101;
		16'b1111010110011110 : data_out =  24'b000000000000010001011110;
		16'b1111010110100000 : data_out =  24'b000000000000010001011111;
		16'b1111010110100010 : data_out =  24'b000000000000010001100000;
		16'b1111010110100100 : data_out =  24'b000000000000010001100001;
		16'b1111010110100110 : data_out =  24'b000000000000010001100011;
		16'b1111010110101000 : data_out =  24'b000000000000010001100100;
		16'b1111010110101010 : data_out =  24'b000000000000010001100101;
		16'b1111010110101101 : data_out =  24'b000000000000010001100110;
		16'b1111010110101111 : data_out =  24'b000000000000010001100111;
		16'b1111010110110001 : data_out =  24'b000000000000010001101000;
		16'b1111010110110011 : data_out =  24'b000000000000010001101001;
		16'b1111010110110101 : data_out =  24'b000000000000010001101010;
		16'b1111010110110111 : data_out =  24'b000000000000010001101100;
		16'b1111010110111001 : data_out =  24'b000000000000010001101101;
		16'b1111010110111011 : data_out =  24'b000000000000010001101110;
		16'b1111010110111101 : data_out =  24'b000000000000010001101111;
		16'b1111010110111111 : data_out =  24'b000000000000010001110000;
		16'b1111010111000001 : data_out =  24'b000000000000010001110001;
		16'b1111010111000011 : data_out =  24'b000000000000010001110010;
		16'b1111010111000101 : data_out =  24'b000000000000010001110011;
		16'b1111010111000111 : data_out =  24'b000000000000010001110101;
		16'b1111010111001001 : data_out =  24'b000000000000010001110110;
		16'b1111010111001011 : data_out =  24'b000000000000010001110111;
		16'b1111010111001101 : data_out =  24'b000000000000010001111000;
		16'b1111010111001111 : data_out =  24'b000000000000010001111001;
		16'b1111010111010001 : data_out =  24'b000000000000010001111010;
		16'b1111010111010011 : data_out =  24'b000000000000010001111011;
		16'b1111010111010101 : data_out =  24'b000000000000010001111101;
		16'b1111010111011000 : data_out =  24'b000000000000010001111110;
		16'b1111010111011010 : data_out =  24'b000000000000010001111111;
		16'b1111010111011100 : data_out =  24'b000000000000010010000000;
		16'b1111010111011110 : data_out =  24'b000000000000010010000001;
		16'b1111010111100000 : data_out =  24'b000000000000010010000010;
		16'b1111010111100010 : data_out =  24'b000000000000010010000100;
		16'b1111010111100100 : data_out =  24'b000000000000010010000101;
		16'b1111010111100110 : data_out =  24'b000000000000010010000110;
		16'b1111010111101000 : data_out =  24'b000000000000010010000111;
		16'b1111010111101010 : data_out =  24'b000000000000010010001000;
		16'b1111010111101100 : data_out =  24'b000000000000010010001001;
		16'b1111010111101110 : data_out =  24'b000000000000010010001011;
		16'b1111010111110000 : data_out =  24'b000000000000010010001100;
		16'b1111010111110010 : data_out =  24'b000000000000010010001101;
		16'b1111010111110100 : data_out =  24'b000000000000010010001110;
		16'b1111010111110110 : data_out =  24'b000000000000010010001111;
		16'b1111010111111000 : data_out =  24'b000000000000010010010000;
		16'b1111010111111010 : data_out =  24'b000000000000010010010010;
		16'b1111010111111100 : data_out =  24'b000000000000010010010011;
		16'b1111010111111110 : data_out =  24'b000000000000010010010100;
		16'b1111011000000001 : data_out =  24'b000000000000010010010101;
		16'b1111011000000011 : data_out =  24'b000000000000010010010110;
		16'b1111011000000101 : data_out =  24'b000000000000010010010111;
		16'b1111011000000111 : data_out =  24'b000000000000010010011001;
		16'b1111011000001001 : data_out =  24'b000000000000010010011010;
		16'b1111011000001011 : data_out =  24'b000000000000010010011011;
		16'b1111011000001101 : data_out =  24'b000000000000010010011100;
		16'b1111011000001111 : data_out =  24'b000000000000010010011101;
		16'b1111011000010001 : data_out =  24'b000000000000010010011110;
		16'b1111011000010011 : data_out =  24'b000000000000010010100000;
		16'b1111011000010101 : data_out =  24'b000000000000010010100001;
		16'b1111011000010111 : data_out =  24'b000000000000010010100010;
		16'b1111011000011001 : data_out =  24'b000000000000010010100011;
		16'b1111011000011011 : data_out =  24'b000000000000010010100100;
		16'b1111011000011101 : data_out =  24'b000000000000010010100110;
		16'b1111011000011111 : data_out =  24'b000000000000010010100111;
		16'b1111011000100001 : data_out =  24'b000000000000010010101000;
		16'b1111011000100011 : data_out =  24'b000000000000010010101001;
		16'b1111011000100101 : data_out =  24'b000000000000010010101010;
		16'b1111011000100111 : data_out =  24'b000000000000010010101100;
		16'b1111011000101001 : data_out =  24'b000000000000010010101101;
		16'b1111011000101100 : data_out =  24'b000000000000010010101110;
		16'b1111011000101110 : data_out =  24'b000000000000010010101111;
		16'b1111011000110000 : data_out =  24'b000000000000010010110000;
		16'b1111011000110010 : data_out =  24'b000000000000010010110010;
		16'b1111011000110100 : data_out =  24'b000000000000010010110011;
		16'b1111011000110110 : data_out =  24'b000000000000010010110100;
		16'b1111011000111000 : data_out =  24'b000000000000010010110101;
		16'b1111011000111010 : data_out =  24'b000000000000010010110110;
		16'b1111011000111100 : data_out =  24'b000000000000010010111000;
		16'b1111011000111110 : data_out =  24'b000000000000010010111001;
		16'b1111011001000000 : data_out =  24'b000000000000010010111010;
		16'b1111011001000010 : data_out =  24'b000000000000010010111011;
		16'b1111011001000100 : data_out =  24'b000000000000010010111100;
		16'b1111011001000110 : data_out =  24'b000000000000010010111110;
		16'b1111011001001000 : data_out =  24'b000000000000010010111111;
		16'b1111011001001010 : data_out =  24'b000000000000010011000000;
		16'b1111011001001100 : data_out =  24'b000000000000010011000001;
		16'b1111011001001110 : data_out =  24'b000000000000010011000010;
		16'b1111011001010000 : data_out =  24'b000000000000010011000100;
		16'b1111011001010010 : data_out =  24'b000000000000010011000101;
		16'b1111011001010100 : data_out =  24'b000000000000010011000110;
		16'b1111011001010111 : data_out =  24'b000000000000010011000111;
		16'b1111011001011001 : data_out =  24'b000000000000010011001001;
		16'b1111011001011011 : data_out =  24'b000000000000010011001010;
		16'b1111011001011101 : data_out =  24'b000000000000010011001011;
		16'b1111011001011111 : data_out =  24'b000000000000010011001100;
		16'b1111011001100001 : data_out =  24'b000000000000010011001101;
		16'b1111011001100011 : data_out =  24'b000000000000010011001111;
		16'b1111011001100101 : data_out =  24'b000000000000010011010000;
		16'b1111011001100111 : data_out =  24'b000000000000010011010001;
		16'b1111011001101001 : data_out =  24'b000000000000010011010010;
		16'b1111011001101011 : data_out =  24'b000000000000010011010100;
		16'b1111011001101101 : data_out =  24'b000000000000010011010101;
		16'b1111011001101111 : data_out =  24'b000000000000010011010110;
		16'b1111011001110001 : data_out =  24'b000000000000010011010111;
		16'b1111011001110011 : data_out =  24'b000000000000010011011001;
		16'b1111011001110101 : data_out =  24'b000000000000010011011010;
		16'b1111011001110111 : data_out =  24'b000000000000010011011011;
		16'b1111011001111001 : data_out =  24'b000000000000010011011100;
		16'b1111011001111011 : data_out =  24'b000000000000010011011110;
		16'b1111011001111101 : data_out =  24'b000000000000010011011111;
		16'b1111011001111111 : data_out =  24'b000000000000010011100000;
		16'b1111011010000010 : data_out =  24'b000000000000010011100001;
		16'b1111011010000100 : data_out =  24'b000000000000010011100011;
		16'b1111011010000110 : data_out =  24'b000000000000010011100100;
		16'b1111011010001000 : data_out =  24'b000000000000010011100101;
		16'b1111011010001010 : data_out =  24'b000000000000010011100110;
		16'b1111011010001100 : data_out =  24'b000000000000010011101000;
		16'b1111011010001110 : data_out =  24'b000000000000010011101001;
		16'b1111011010010000 : data_out =  24'b000000000000010011101010;
		16'b1111011010010010 : data_out =  24'b000000000000010011101011;
		16'b1111011010010100 : data_out =  24'b000000000000010011101101;
		16'b1111011010010110 : data_out =  24'b000000000000010011101110;
		16'b1111011010011000 : data_out =  24'b000000000000010011101111;
		16'b1111011010011010 : data_out =  24'b000000000000010011110000;
		16'b1111011010011100 : data_out =  24'b000000000000010011110010;
		16'b1111011010011110 : data_out =  24'b000000000000010011110011;
		16'b1111011010100000 : data_out =  24'b000000000000010011110100;
		16'b1111011010100010 : data_out =  24'b000000000000010011110101;
		16'b1111011010100100 : data_out =  24'b000000000000010011110111;
		16'b1111011010100110 : data_out =  24'b000000000000010011111000;
		16'b1111011010101000 : data_out =  24'b000000000000010011111001;
		16'b1111011010101010 : data_out =  24'b000000000000010011111011;
		16'b1111011010101101 : data_out =  24'b000000000000010011111100;
		16'b1111011010101111 : data_out =  24'b000000000000010011111101;
		16'b1111011010110001 : data_out =  24'b000000000000010011111110;
		16'b1111011010110011 : data_out =  24'b000000000000010100000000;
		16'b1111011010110101 : data_out =  24'b000000000000010100000001;
		16'b1111011010110111 : data_out =  24'b000000000000010100000010;
		16'b1111011010111001 : data_out =  24'b000000000000010100000100;
		16'b1111011010111011 : data_out =  24'b000000000000010100000101;
		16'b1111011010111101 : data_out =  24'b000000000000010100000110;
		16'b1111011010111111 : data_out =  24'b000000000000010100000111;
		16'b1111011011000001 : data_out =  24'b000000000000010100001001;
		16'b1111011011000011 : data_out =  24'b000000000000010100001010;
		16'b1111011011000101 : data_out =  24'b000000000000010100001011;
		16'b1111011011000111 : data_out =  24'b000000000000010100001101;
		16'b1111011011001001 : data_out =  24'b000000000000010100001110;
		16'b1111011011001011 : data_out =  24'b000000000000010100001111;
		16'b1111011011001101 : data_out =  24'b000000000000010100010000;
		16'b1111011011001111 : data_out =  24'b000000000000010100010010;
		16'b1111011011010001 : data_out =  24'b000000000000010100010011;
		16'b1111011011010011 : data_out =  24'b000000000000010100010100;
		16'b1111011011010101 : data_out =  24'b000000000000010100010110;
		16'b1111011011011000 : data_out =  24'b000000000000010100010111;
		16'b1111011011011010 : data_out =  24'b000000000000010100011000;
		16'b1111011011011100 : data_out =  24'b000000000000010100011010;
		16'b1111011011011110 : data_out =  24'b000000000000010100011011;
		16'b1111011011100000 : data_out =  24'b000000000000010100011100;
		16'b1111011011100010 : data_out =  24'b000000000000010100011101;
		16'b1111011011100100 : data_out =  24'b000000000000010100011111;
		16'b1111011011100110 : data_out =  24'b000000000000010100100000;
		16'b1111011011101000 : data_out =  24'b000000000000010100100001;
		16'b1111011011101010 : data_out =  24'b000000000000010100100011;
		16'b1111011011101100 : data_out =  24'b000000000000010100100100;
		16'b1111011011101110 : data_out =  24'b000000000000010100100101;
		16'b1111011011110000 : data_out =  24'b000000000000010100100111;
		16'b1111011011110010 : data_out =  24'b000000000000010100101000;
		16'b1111011011110100 : data_out =  24'b000000000000010100101001;
		16'b1111011011110110 : data_out =  24'b000000000000010100101011;
		16'b1111011011111000 : data_out =  24'b000000000000010100101100;
		16'b1111011011111010 : data_out =  24'b000000000000010100101101;
		16'b1111011011111100 : data_out =  24'b000000000000010100101111;
		16'b1111011011111110 : data_out =  24'b000000000000010100110000;
		16'b1111011100000001 : data_out =  24'b000000000000010100110001;
		16'b1111011100000011 : data_out =  24'b000000000000010100110011;
		16'b1111011100000101 : data_out =  24'b000000000000010100110100;
		16'b1111011100000111 : data_out =  24'b000000000000010100110101;
		16'b1111011100001001 : data_out =  24'b000000000000010100110111;
		16'b1111011100001011 : data_out =  24'b000000000000010100111000;
		16'b1111011100001101 : data_out =  24'b000000000000010100111001;
		16'b1111011100001111 : data_out =  24'b000000000000010100111011;
		16'b1111011100010001 : data_out =  24'b000000000000010100111100;
		16'b1111011100010011 : data_out =  24'b000000000000010100111101;
		16'b1111011100010101 : data_out =  24'b000000000000010100111111;
		16'b1111011100010111 : data_out =  24'b000000000000010101000000;
		16'b1111011100011001 : data_out =  24'b000000000000010101000001;
		16'b1111011100011011 : data_out =  24'b000000000000010101000011;
		16'b1111011100011101 : data_out =  24'b000000000000010101000100;
		16'b1111011100011111 : data_out =  24'b000000000000010101000101;
		16'b1111011100100001 : data_out =  24'b000000000000010101000111;
		16'b1111011100100011 : data_out =  24'b000000000000010101001000;
		16'b1111011100100101 : data_out =  24'b000000000000010101001001;
		16'b1111011100100111 : data_out =  24'b000000000000010101001011;
		16'b1111011100101001 : data_out =  24'b000000000000010101001100;
		16'b1111011100101100 : data_out =  24'b000000000000010101001101;
		16'b1111011100101110 : data_out =  24'b000000000000010101001111;
		16'b1111011100110000 : data_out =  24'b000000000000010101010000;
		16'b1111011100110010 : data_out =  24'b000000000000010101010010;
		16'b1111011100110100 : data_out =  24'b000000000000010101010011;
		16'b1111011100110110 : data_out =  24'b000000000000010101010100;
		16'b1111011100111000 : data_out =  24'b000000000000010101010110;
		16'b1111011100111010 : data_out =  24'b000000000000010101010111;
		16'b1111011100111100 : data_out =  24'b000000000000010101011000;
		16'b1111011100111110 : data_out =  24'b000000000000010101011010;
		16'b1111011101000000 : data_out =  24'b000000000000010101011011;
		16'b1111011101000010 : data_out =  24'b000000000000010101011101;
		16'b1111011101000100 : data_out =  24'b000000000000010101011110;
		16'b1111011101000110 : data_out =  24'b000000000000010101011111;
		16'b1111011101001000 : data_out =  24'b000000000000010101100001;
		16'b1111011101001010 : data_out =  24'b000000000000010101100010;
		16'b1111011101001100 : data_out =  24'b000000000000010101100011;
		16'b1111011101001110 : data_out =  24'b000000000000010101100101;
		16'b1111011101010000 : data_out =  24'b000000000000010101100110;
		16'b1111011101010010 : data_out =  24'b000000000000010101101000;
		16'b1111011101010100 : data_out =  24'b000000000000010101101001;
		16'b1111011101010111 : data_out =  24'b000000000000010101101010;
		16'b1111011101011001 : data_out =  24'b000000000000010101101100;
		16'b1111011101011011 : data_out =  24'b000000000000010101101101;
		16'b1111011101011101 : data_out =  24'b000000000000010101101110;
		16'b1111011101011111 : data_out =  24'b000000000000010101110000;
		16'b1111011101100001 : data_out =  24'b000000000000010101110001;
		16'b1111011101100011 : data_out =  24'b000000000000010101110011;
		16'b1111011101100101 : data_out =  24'b000000000000010101110100;
		16'b1111011101100111 : data_out =  24'b000000000000010101110101;
		16'b1111011101101001 : data_out =  24'b000000000000010101110111;
		16'b1111011101101011 : data_out =  24'b000000000000010101111000;
		16'b1111011101101101 : data_out =  24'b000000000000010101111010;
		16'b1111011101101111 : data_out =  24'b000000000000010101111011;
		16'b1111011101110001 : data_out =  24'b000000000000010101111100;
		16'b1111011101110011 : data_out =  24'b000000000000010101111110;
		16'b1111011101110101 : data_out =  24'b000000000000010101111111;
		16'b1111011101110111 : data_out =  24'b000000000000010110000001;
		16'b1111011101111001 : data_out =  24'b000000000000010110000010;
		16'b1111011101111011 : data_out =  24'b000000000000010110000100;
		16'b1111011101111101 : data_out =  24'b000000000000010110000101;
		16'b1111011101111111 : data_out =  24'b000000000000010110000110;
		16'b1111011110000010 : data_out =  24'b000000000000010110001000;
		16'b1111011110000100 : data_out =  24'b000000000000010110001001;
		16'b1111011110000110 : data_out =  24'b000000000000010110001011;
		16'b1111011110001000 : data_out =  24'b000000000000010110001100;
		16'b1111011110001010 : data_out =  24'b000000000000010110001101;
		16'b1111011110001100 : data_out =  24'b000000000000010110001111;
		16'b1111011110001110 : data_out =  24'b000000000000010110010000;
		16'b1111011110010000 : data_out =  24'b000000000000010110010010;
		16'b1111011110010010 : data_out =  24'b000000000000010110010011;
		16'b1111011110010100 : data_out =  24'b000000000000010110010101;
		16'b1111011110010110 : data_out =  24'b000000000000010110010110;
		16'b1111011110011000 : data_out =  24'b000000000000010110010111;
		16'b1111011110011010 : data_out =  24'b000000000000010110011001;
		16'b1111011110011100 : data_out =  24'b000000000000010110011010;
		16'b1111011110011110 : data_out =  24'b000000000000010110011100;
		16'b1111011110100000 : data_out =  24'b000000000000010110011101;
		16'b1111011110100010 : data_out =  24'b000000000000010110011111;
		16'b1111011110100100 : data_out =  24'b000000000000010110100000;
		16'b1111011110100110 : data_out =  24'b000000000000010110100001;
		16'b1111011110101000 : data_out =  24'b000000000000010110100011;
		16'b1111011110101010 : data_out =  24'b000000000000010110100100;
		16'b1111011110101101 : data_out =  24'b000000000000010110100110;
		16'b1111011110101111 : data_out =  24'b000000000000010110100111;
		16'b1111011110110001 : data_out =  24'b000000000000010110101001;
		16'b1111011110110011 : data_out =  24'b000000000000010110101010;
		16'b1111011110110101 : data_out =  24'b000000000000010110101100;
		16'b1111011110110111 : data_out =  24'b000000000000010110101101;
		16'b1111011110111001 : data_out =  24'b000000000000010110101111;
		16'b1111011110111011 : data_out =  24'b000000000000010110110000;
		16'b1111011110111101 : data_out =  24'b000000000000010110110001;
		16'b1111011110111111 : data_out =  24'b000000000000010110110011;
		16'b1111011111000001 : data_out =  24'b000000000000010110110100;
		16'b1111011111000011 : data_out =  24'b000000000000010110110110;
		16'b1111011111000101 : data_out =  24'b000000000000010110110111;
		16'b1111011111000111 : data_out =  24'b000000000000010110111001;
		16'b1111011111001001 : data_out =  24'b000000000000010110111010;
		16'b1111011111001011 : data_out =  24'b000000000000010110111100;
		16'b1111011111001101 : data_out =  24'b000000000000010110111101;
		16'b1111011111001111 : data_out =  24'b000000000000010110111111;
		16'b1111011111010001 : data_out =  24'b000000000000010111000000;
		16'b1111011111010011 : data_out =  24'b000000000000010111000010;
		16'b1111011111010101 : data_out =  24'b000000000000010111000011;
		16'b1111011111011000 : data_out =  24'b000000000000010111000100;
		16'b1111011111011010 : data_out =  24'b000000000000010111000110;
		16'b1111011111011100 : data_out =  24'b000000000000010111000111;
		16'b1111011111011110 : data_out =  24'b000000000000010111001001;
		16'b1111011111100000 : data_out =  24'b000000000000010111001010;
		16'b1111011111100010 : data_out =  24'b000000000000010111001100;
		16'b1111011111100100 : data_out =  24'b000000000000010111001101;
		16'b1111011111100110 : data_out =  24'b000000000000010111001111;
		16'b1111011111101000 : data_out =  24'b000000000000010111010000;
		16'b1111011111101010 : data_out =  24'b000000000000010111010010;
		16'b1111011111101100 : data_out =  24'b000000000000010111010011;
		16'b1111011111101110 : data_out =  24'b000000000000010111010101;
		16'b1111011111110000 : data_out =  24'b000000000000010111010110;
		16'b1111011111110010 : data_out =  24'b000000000000010111011000;
		16'b1111011111110100 : data_out =  24'b000000000000010111011001;
		16'b1111011111110110 : data_out =  24'b000000000000010111011011;
		16'b1111011111111000 : data_out =  24'b000000000000010111011100;
		16'b1111011111111010 : data_out =  24'b000000000000010111011110;
		16'b1111011111111100 : data_out =  24'b000000000000010111011111;
		16'b1111011111111110 : data_out =  24'b000000000000010111100001;
		16'b1111100000000001 : data_out =  24'b000000000000010111100010;
		16'b1111100000000011 : data_out =  24'b000000000000010111100100;
		16'b1111100000000101 : data_out =  24'b000000000000010111100101;
		16'b1111100000000111 : data_out =  24'b000000000000010111100111;
		16'b1111100000001001 : data_out =  24'b000000000000010111101000;
		16'b1111100000001011 : data_out =  24'b000000000000010111101010;
		16'b1111100000001101 : data_out =  24'b000000000000010111101011;
		16'b1111100000001111 : data_out =  24'b000000000000010111101101;
		16'b1111100000010001 : data_out =  24'b000000000000010111101110;
		16'b1111100000010011 : data_out =  24'b000000000000010111110000;
		16'b1111100000010101 : data_out =  24'b000000000000010111110001;
		16'b1111100000010111 : data_out =  24'b000000000000010111110011;
		16'b1111100000011001 : data_out =  24'b000000000000010111110101;
		16'b1111100000011011 : data_out =  24'b000000000000010111110110;
		16'b1111100000011101 : data_out =  24'b000000000000010111111000;
		16'b1111100000011111 : data_out =  24'b000000000000010111111001;
		16'b1111100000100001 : data_out =  24'b000000000000010111111011;
		16'b1111100000100011 : data_out =  24'b000000000000010111111100;
		16'b1111100000100101 : data_out =  24'b000000000000010111111110;
		16'b1111100000100111 : data_out =  24'b000000000000010111111111;
		16'b1111100000101001 : data_out =  24'b000000000000011000000001;
		16'b1111100000101100 : data_out =  24'b000000000000011000000010;
		16'b1111100000101110 : data_out =  24'b000000000000011000000100;
		16'b1111100000110000 : data_out =  24'b000000000000011000000101;
		16'b1111100000110010 : data_out =  24'b000000000000011000000111;
		16'b1111100000110100 : data_out =  24'b000000000000011000001000;
		16'b1111100000110110 : data_out =  24'b000000000000011000001010;
		16'b1111100000111000 : data_out =  24'b000000000000011000001100;
		16'b1111100000111010 : data_out =  24'b000000000000011000001101;
		16'b1111100000111100 : data_out =  24'b000000000000011000001111;
		16'b1111100000111110 : data_out =  24'b000000000000011000010000;
		16'b1111100001000000 : data_out =  24'b000000000000011000010010;
		16'b1111100001000010 : data_out =  24'b000000000000011000010011;
		16'b1111100001000100 : data_out =  24'b000000000000011000010101;
		16'b1111100001000110 : data_out =  24'b000000000000011000010110;
		16'b1111100001001000 : data_out =  24'b000000000000011000011000;
		16'b1111100001001010 : data_out =  24'b000000000000011000011010;
		16'b1111100001001100 : data_out =  24'b000000000000011000011011;
		16'b1111100001001110 : data_out =  24'b000000000000011000011101;
		16'b1111100001010000 : data_out =  24'b000000000000011000011110;
		16'b1111100001010010 : data_out =  24'b000000000000011000100000;
		16'b1111100001010100 : data_out =  24'b000000000000011000100001;
		16'b1111100001010111 : data_out =  24'b000000000000011000100011;
		16'b1111100001011001 : data_out =  24'b000000000000011000100101;
		16'b1111100001011011 : data_out =  24'b000000000000011000100110;
		16'b1111100001011101 : data_out =  24'b000000000000011000101000;
		16'b1111100001011111 : data_out =  24'b000000000000011000101001;
		16'b1111100001100001 : data_out =  24'b000000000000011000101011;
		16'b1111100001100011 : data_out =  24'b000000000000011000101100;
		16'b1111100001100101 : data_out =  24'b000000000000011000101110;
		16'b1111100001100111 : data_out =  24'b000000000000011000110000;
		16'b1111100001101001 : data_out =  24'b000000000000011000110001;
		16'b1111100001101011 : data_out =  24'b000000000000011000110011;
		16'b1111100001101101 : data_out =  24'b000000000000011000110100;
		16'b1111100001101111 : data_out =  24'b000000000000011000110110;
		16'b1111100001110001 : data_out =  24'b000000000000011000111000;
		16'b1111100001110011 : data_out =  24'b000000000000011000111001;
		16'b1111100001110101 : data_out =  24'b000000000000011000111011;
		16'b1111100001110111 : data_out =  24'b000000000000011000111100;
		16'b1111100001111001 : data_out =  24'b000000000000011000111110;
		16'b1111100001111011 : data_out =  24'b000000000000011001000000;
		16'b1111100001111101 : data_out =  24'b000000000000011001000001;
		16'b1111100001111111 : data_out =  24'b000000000000011001000011;
		16'b1111100010000010 : data_out =  24'b000000000000011001000100;
		16'b1111100010000100 : data_out =  24'b000000000000011001000110;
		16'b1111100010000110 : data_out =  24'b000000000000011001001000;
		16'b1111100010001000 : data_out =  24'b000000000000011001001001;
		16'b1111100010001010 : data_out =  24'b000000000000011001001011;
		16'b1111100010001100 : data_out =  24'b000000000000011001001100;
		16'b1111100010001110 : data_out =  24'b000000000000011001001110;
		16'b1111100010010000 : data_out =  24'b000000000000011001010000;
		16'b1111100010010010 : data_out =  24'b000000000000011001010001;
		16'b1111100010010100 : data_out =  24'b000000000000011001010011;
		16'b1111100010010110 : data_out =  24'b000000000000011001010100;
		16'b1111100010011000 : data_out =  24'b000000000000011001010110;
		16'b1111100010011010 : data_out =  24'b000000000000011001011000;
		16'b1111100010011100 : data_out =  24'b000000000000011001011001;
		16'b1111100010011110 : data_out =  24'b000000000000011001011011;
		16'b1111100010100000 : data_out =  24'b000000000000011001011101;
		16'b1111100010100010 : data_out =  24'b000000000000011001011110;
		16'b1111100010100100 : data_out =  24'b000000000000011001100000;
		16'b1111100010100110 : data_out =  24'b000000000000011001100001;
		16'b1111100010101000 : data_out =  24'b000000000000011001100011;
		16'b1111100010101010 : data_out =  24'b000000000000011001100101;
		16'b1111100010101101 : data_out =  24'b000000000000011001100110;
		16'b1111100010101111 : data_out =  24'b000000000000011001101000;
		16'b1111100010110001 : data_out =  24'b000000000000011001101010;
		16'b1111100010110011 : data_out =  24'b000000000000011001101011;
		16'b1111100010110101 : data_out =  24'b000000000000011001101101;
		16'b1111100010110111 : data_out =  24'b000000000000011001101111;
		16'b1111100010111001 : data_out =  24'b000000000000011001110000;
		16'b1111100010111011 : data_out =  24'b000000000000011001110010;
		16'b1111100010111101 : data_out =  24'b000000000000011001110100;
		16'b1111100010111111 : data_out =  24'b000000000000011001110101;
		16'b1111100011000001 : data_out =  24'b000000000000011001110111;
		16'b1111100011000011 : data_out =  24'b000000000000011001111001;
		16'b1111100011000101 : data_out =  24'b000000000000011001111010;
		16'b1111100011000111 : data_out =  24'b000000000000011001111100;
		16'b1111100011001001 : data_out =  24'b000000000000011001111101;
		16'b1111100011001011 : data_out =  24'b000000000000011001111111;
		16'b1111100011001101 : data_out =  24'b000000000000011010000001;
		16'b1111100011001111 : data_out =  24'b000000000000011010000010;
		16'b1111100011010001 : data_out =  24'b000000000000011010000100;
		16'b1111100011010011 : data_out =  24'b000000000000011010000110;
		16'b1111100011010101 : data_out =  24'b000000000000011010000111;
		16'b1111100011011000 : data_out =  24'b000000000000011010001001;
		16'b1111100011011010 : data_out =  24'b000000000000011010001011;
		16'b1111100011011100 : data_out =  24'b000000000000011010001101;
		16'b1111100011011110 : data_out =  24'b000000000000011010001110;
		16'b1111100011100000 : data_out =  24'b000000000000011010010000;
		16'b1111100011100010 : data_out =  24'b000000000000011010010010;
		16'b1111100011100100 : data_out =  24'b000000000000011010010011;
		16'b1111100011100110 : data_out =  24'b000000000000011010010101;
		16'b1111100011101000 : data_out =  24'b000000000000011010010111;
		16'b1111100011101010 : data_out =  24'b000000000000011010011000;
		16'b1111100011101100 : data_out =  24'b000000000000011010011010;
		16'b1111100011101110 : data_out =  24'b000000000000011010011100;
		16'b1111100011110000 : data_out =  24'b000000000000011010011101;
		16'b1111100011110010 : data_out =  24'b000000000000011010011111;
		16'b1111100011110100 : data_out =  24'b000000000000011010100001;
		16'b1111100011110110 : data_out =  24'b000000000000011010100010;
		16'b1111100011111000 : data_out =  24'b000000000000011010100100;
		16'b1111100011111010 : data_out =  24'b000000000000011010100110;
		16'b1111100011111100 : data_out =  24'b000000000000011010101000;
		16'b1111100011111110 : data_out =  24'b000000000000011010101001;
		16'b1111100100000001 : data_out =  24'b000000000000011010101011;
		16'b1111100100000011 : data_out =  24'b000000000000011010101101;
		16'b1111100100000101 : data_out =  24'b000000000000011010101110;
		16'b1111100100000111 : data_out =  24'b000000000000011010110000;
		16'b1111100100001001 : data_out =  24'b000000000000011010110010;
		16'b1111100100001011 : data_out =  24'b000000000000011010110100;
		16'b1111100100001101 : data_out =  24'b000000000000011010110101;
		16'b1111100100001111 : data_out =  24'b000000000000011010110111;
		16'b1111100100010001 : data_out =  24'b000000000000011010111001;
		16'b1111100100010011 : data_out =  24'b000000000000011010111010;
		16'b1111100100010101 : data_out =  24'b000000000000011010111100;
		16'b1111100100010111 : data_out =  24'b000000000000011010111110;
		16'b1111100100011001 : data_out =  24'b000000000000011011000000;
		16'b1111100100011011 : data_out =  24'b000000000000011011000001;
		16'b1111100100011101 : data_out =  24'b000000000000011011000011;
		16'b1111100100011111 : data_out =  24'b000000000000011011000101;
		16'b1111100100100001 : data_out =  24'b000000000000011011000111;
		16'b1111100100100011 : data_out =  24'b000000000000011011001000;
		16'b1111100100100101 : data_out =  24'b000000000000011011001010;
		16'b1111100100100111 : data_out =  24'b000000000000011011001100;
		16'b1111100100101001 : data_out =  24'b000000000000011011001101;
		16'b1111100100101100 : data_out =  24'b000000000000011011001111;
		16'b1111100100101110 : data_out =  24'b000000000000011011010001;
		16'b1111100100110000 : data_out =  24'b000000000000011011010011;
		16'b1111100100110010 : data_out =  24'b000000000000011011010100;
		16'b1111100100110100 : data_out =  24'b000000000000011011010110;
		16'b1111100100110110 : data_out =  24'b000000000000011011011000;
		16'b1111100100111000 : data_out =  24'b000000000000011011011010;
		16'b1111100100111010 : data_out =  24'b000000000000011011011011;
		16'b1111100100111100 : data_out =  24'b000000000000011011011101;
		16'b1111100100111110 : data_out =  24'b000000000000011011011111;
		16'b1111100101000000 : data_out =  24'b000000000000011011100001;
		16'b1111100101000010 : data_out =  24'b000000000000011011100010;
		16'b1111100101000100 : data_out =  24'b000000000000011011100100;
		16'b1111100101000110 : data_out =  24'b000000000000011011100110;
		16'b1111100101001000 : data_out =  24'b000000000000011011101000;
		16'b1111100101001010 : data_out =  24'b000000000000011011101010;
		16'b1111100101001100 : data_out =  24'b000000000000011011101011;
		16'b1111100101001110 : data_out =  24'b000000000000011011101101;
		16'b1111100101010000 : data_out =  24'b000000000000011011101111;
		16'b1111100101010010 : data_out =  24'b000000000000011011110001;
		16'b1111100101010100 : data_out =  24'b000000000000011011110010;
		16'b1111100101010111 : data_out =  24'b000000000000011011110100;
		16'b1111100101011001 : data_out =  24'b000000000000011011110110;
		16'b1111100101011011 : data_out =  24'b000000000000011011111000;
		16'b1111100101011101 : data_out =  24'b000000000000011011111010;
		16'b1111100101011111 : data_out =  24'b000000000000011011111011;
		16'b1111100101100001 : data_out =  24'b000000000000011011111101;
		16'b1111100101100011 : data_out =  24'b000000000000011011111111;
		16'b1111100101100101 : data_out =  24'b000000000000011100000001;
		16'b1111100101100111 : data_out =  24'b000000000000011100000011;
		16'b1111100101101001 : data_out =  24'b000000000000011100000100;
		16'b1111100101101011 : data_out =  24'b000000000000011100000110;
		16'b1111100101101101 : data_out =  24'b000000000000011100001000;
		16'b1111100101101111 : data_out =  24'b000000000000011100001010;
		16'b1111100101110001 : data_out =  24'b000000000000011100001100;
		16'b1111100101110011 : data_out =  24'b000000000000011100001101;
		16'b1111100101110101 : data_out =  24'b000000000000011100001111;
		16'b1111100101110111 : data_out =  24'b000000000000011100010001;
		16'b1111100101111001 : data_out =  24'b000000000000011100010011;
		16'b1111100101111011 : data_out =  24'b000000000000011100010101;
		16'b1111100101111101 : data_out =  24'b000000000000011100010110;
		16'b1111100101111111 : data_out =  24'b000000000000011100011000;
		16'b1111100110000010 : data_out =  24'b000000000000011100011010;
		16'b1111100110000100 : data_out =  24'b000000000000011100011100;
		16'b1111100110000110 : data_out =  24'b000000000000011100011110;
		16'b1111100110001000 : data_out =  24'b000000000000011100011111;
		16'b1111100110001010 : data_out =  24'b000000000000011100100001;
		16'b1111100110001100 : data_out =  24'b000000000000011100100011;
		16'b1111100110001110 : data_out =  24'b000000000000011100100101;
		16'b1111100110010000 : data_out =  24'b000000000000011100100111;
		16'b1111100110010010 : data_out =  24'b000000000000011100101001;
		16'b1111100110010100 : data_out =  24'b000000000000011100101010;
		16'b1111100110010110 : data_out =  24'b000000000000011100101100;
		16'b1111100110011000 : data_out =  24'b000000000000011100101110;
		16'b1111100110011010 : data_out =  24'b000000000000011100110000;
		16'b1111100110011100 : data_out =  24'b000000000000011100110010;
		16'b1111100110011110 : data_out =  24'b000000000000011100110100;
		16'b1111100110100000 : data_out =  24'b000000000000011100110101;
		16'b1111100110100010 : data_out =  24'b000000000000011100110111;
		16'b1111100110100100 : data_out =  24'b000000000000011100111001;
		16'b1111100110100110 : data_out =  24'b000000000000011100111011;
		16'b1111100110101000 : data_out =  24'b000000000000011100111101;
		16'b1111100110101010 : data_out =  24'b000000000000011100111111;
		16'b1111100110101101 : data_out =  24'b000000000000011101000001;
		16'b1111100110101111 : data_out =  24'b000000000000011101000010;
		16'b1111100110110001 : data_out =  24'b000000000000011101000100;
		16'b1111100110110011 : data_out =  24'b000000000000011101000110;
		16'b1111100110110101 : data_out =  24'b000000000000011101001000;
		16'b1111100110110111 : data_out =  24'b000000000000011101001010;
		16'b1111100110111001 : data_out =  24'b000000000000011101001100;
		16'b1111100110111011 : data_out =  24'b000000000000011101001110;
		16'b1111100110111101 : data_out =  24'b000000000000011101010000;
		16'b1111100110111111 : data_out =  24'b000000000000011101010001;
		16'b1111100111000001 : data_out =  24'b000000000000011101010011;
		16'b1111100111000011 : data_out =  24'b000000000000011101010101;
		16'b1111100111000101 : data_out =  24'b000000000000011101010111;
		16'b1111100111000111 : data_out =  24'b000000000000011101011001;
		16'b1111100111001001 : data_out =  24'b000000000000011101011011;
		16'b1111100111001011 : data_out =  24'b000000000000011101011101;
		16'b1111100111001101 : data_out =  24'b000000000000011101011111;
		16'b1111100111001111 : data_out =  24'b000000000000011101100000;
		16'b1111100111010001 : data_out =  24'b000000000000011101100010;
		16'b1111100111010011 : data_out =  24'b000000000000011101100100;
		16'b1111100111010101 : data_out =  24'b000000000000011101100110;
		16'b1111100111011000 : data_out =  24'b000000000000011101101000;
		16'b1111100111011010 : data_out =  24'b000000000000011101101010;
		16'b1111100111011100 : data_out =  24'b000000000000011101101100;
		16'b1111100111011110 : data_out =  24'b000000000000011101101110;
		16'b1111100111100000 : data_out =  24'b000000000000011101110000;
		16'b1111100111100010 : data_out =  24'b000000000000011101110010;
		16'b1111100111100100 : data_out =  24'b000000000000011101110011;
		16'b1111100111100110 : data_out =  24'b000000000000011101110101;
		16'b1111100111101000 : data_out =  24'b000000000000011101110111;
		16'b1111100111101010 : data_out =  24'b000000000000011101111001;
		16'b1111100111101100 : data_out =  24'b000000000000011101111011;
		16'b1111100111101110 : data_out =  24'b000000000000011101111101;
		16'b1111100111110000 : data_out =  24'b000000000000011101111111;
		16'b1111100111110010 : data_out =  24'b000000000000011110000001;
		16'b1111100111110100 : data_out =  24'b000000000000011110000011;
		16'b1111100111110110 : data_out =  24'b000000000000011110000101;
		16'b1111100111111000 : data_out =  24'b000000000000011110000111;
		16'b1111100111111010 : data_out =  24'b000000000000011110001001;
		16'b1111100111111100 : data_out =  24'b000000000000011110001010;
		16'b1111100111111110 : data_out =  24'b000000000000011110001100;
		16'b1111101000000001 : data_out =  24'b000000000000011110001110;
		16'b1111101000000011 : data_out =  24'b000000000000011110010000;
		16'b1111101000000101 : data_out =  24'b000000000000011110010010;
		16'b1111101000000111 : data_out =  24'b000000000000011110010100;
		16'b1111101000001001 : data_out =  24'b000000000000011110010110;
		16'b1111101000001011 : data_out =  24'b000000000000011110011000;
		16'b1111101000001101 : data_out =  24'b000000000000011110011010;
		16'b1111101000001111 : data_out =  24'b000000000000011110011100;
		16'b1111101000010001 : data_out =  24'b000000000000011110011110;
		16'b1111101000010011 : data_out =  24'b000000000000011110100000;
		16'b1111101000010101 : data_out =  24'b000000000000011110100010;
		16'b1111101000010111 : data_out =  24'b000000000000011110100100;
		16'b1111101000011001 : data_out =  24'b000000000000011110100110;
		16'b1111101000011011 : data_out =  24'b000000000000011110101000;
		16'b1111101000011101 : data_out =  24'b000000000000011110101010;
		16'b1111101000011111 : data_out =  24'b000000000000011110101100;
		16'b1111101000100001 : data_out =  24'b000000000000011110101110;
		16'b1111101000100011 : data_out =  24'b000000000000011110101111;
		16'b1111101000100101 : data_out =  24'b000000000000011110110001;
		16'b1111101000100111 : data_out =  24'b000000000000011110110011;
		16'b1111101000101001 : data_out =  24'b000000000000011110110101;
		16'b1111101000101100 : data_out =  24'b000000000000011110110111;
		16'b1111101000101110 : data_out =  24'b000000000000011110111001;
		16'b1111101000110000 : data_out =  24'b000000000000011110111011;
		16'b1111101000110010 : data_out =  24'b000000000000011110111101;
		16'b1111101000110100 : data_out =  24'b000000000000011110111111;
		16'b1111101000110110 : data_out =  24'b000000000000011111000001;
		16'b1111101000111000 : data_out =  24'b000000000000011111000011;
		16'b1111101000111010 : data_out =  24'b000000000000011111000101;
		16'b1111101000111100 : data_out =  24'b000000000000011111000111;
		16'b1111101000111110 : data_out =  24'b000000000000011111001001;
		16'b1111101001000000 : data_out =  24'b000000000000011111001011;
		16'b1111101001000010 : data_out =  24'b000000000000011111001101;
		16'b1111101001000100 : data_out =  24'b000000000000011111001111;
		16'b1111101001000110 : data_out =  24'b000000000000011111010001;
		16'b1111101001001000 : data_out =  24'b000000000000011111010011;
		16'b1111101001001010 : data_out =  24'b000000000000011111010101;
		16'b1111101001001100 : data_out =  24'b000000000000011111010111;
		16'b1111101001001110 : data_out =  24'b000000000000011111011001;
		16'b1111101001010000 : data_out =  24'b000000000000011111011011;
		16'b1111101001010010 : data_out =  24'b000000000000011111011101;
		16'b1111101001010100 : data_out =  24'b000000000000011111011111;
		16'b1111101001010111 : data_out =  24'b000000000000011111100001;
		16'b1111101001011001 : data_out =  24'b000000000000011111100011;
		16'b1111101001011011 : data_out =  24'b000000000000011111100101;
		16'b1111101001011101 : data_out =  24'b000000000000011111100111;
		16'b1111101001011111 : data_out =  24'b000000000000011111101001;
		16'b1111101001100001 : data_out =  24'b000000000000011111101011;
		16'b1111101001100011 : data_out =  24'b000000000000011111101101;
		16'b1111101001100101 : data_out =  24'b000000000000011111101111;
		16'b1111101001100111 : data_out =  24'b000000000000011111110010;
		16'b1111101001101001 : data_out =  24'b000000000000011111110100;
		16'b1111101001101011 : data_out =  24'b000000000000011111110110;
		16'b1111101001101101 : data_out =  24'b000000000000011111111000;
		16'b1111101001101111 : data_out =  24'b000000000000011111111010;
		16'b1111101001110001 : data_out =  24'b000000000000011111111100;
		16'b1111101001110011 : data_out =  24'b000000000000011111111110;
		16'b1111101001110101 : data_out =  24'b000000000000100000000000;
		16'b1111101001110111 : data_out =  24'b000000000000100000000010;
		16'b1111101001111001 : data_out =  24'b000000000000100000000100;
		16'b1111101001111011 : data_out =  24'b000000000000100000000110;
		16'b1111101001111101 : data_out =  24'b000000000000100000001000;
		16'b1111101001111111 : data_out =  24'b000000000000100000001010;
		16'b1111101010000010 : data_out =  24'b000000000000100000001100;
		16'b1111101010000100 : data_out =  24'b000000000000100000001110;
		16'b1111101010000110 : data_out =  24'b000000000000100000010000;
		16'b1111101010001000 : data_out =  24'b000000000000100000010010;
		16'b1111101010001010 : data_out =  24'b000000000000100000010100;
		16'b1111101010001100 : data_out =  24'b000000000000100000010110;
		16'b1111101010001110 : data_out =  24'b000000000000100000011001;
		16'b1111101010010000 : data_out =  24'b000000000000100000011011;
		16'b1111101010010010 : data_out =  24'b000000000000100000011101;
		16'b1111101010010100 : data_out =  24'b000000000000100000011111;
		16'b1111101010010110 : data_out =  24'b000000000000100000100001;
		16'b1111101010011000 : data_out =  24'b000000000000100000100011;
		16'b1111101010011010 : data_out =  24'b000000000000100000100101;
		16'b1111101010011100 : data_out =  24'b000000000000100000100111;
		16'b1111101010011110 : data_out =  24'b000000000000100000101001;
		16'b1111101010100000 : data_out =  24'b000000000000100000101011;
		16'b1111101010100010 : data_out =  24'b000000000000100000101101;
		16'b1111101010100100 : data_out =  24'b000000000000100000101111;
		16'b1111101010100110 : data_out =  24'b000000000000100000110010;
		16'b1111101010101000 : data_out =  24'b000000000000100000110100;
		16'b1111101010101010 : data_out =  24'b000000000000100000110110;
		16'b1111101010101101 : data_out =  24'b000000000000100000111000;
		16'b1111101010101111 : data_out =  24'b000000000000100000111010;
		16'b1111101010110001 : data_out =  24'b000000000000100000111100;
		16'b1111101010110011 : data_out =  24'b000000000000100000111110;
		16'b1111101010110101 : data_out =  24'b000000000000100001000000;
		16'b1111101010110111 : data_out =  24'b000000000000100001000010;
		16'b1111101010111001 : data_out =  24'b000000000000100001000101;
		16'b1111101010111011 : data_out =  24'b000000000000100001000111;
		16'b1111101010111101 : data_out =  24'b000000000000100001001001;
		16'b1111101010111111 : data_out =  24'b000000000000100001001011;
		16'b1111101011000001 : data_out =  24'b000000000000100001001101;
		16'b1111101011000011 : data_out =  24'b000000000000100001001111;
		16'b1111101011000101 : data_out =  24'b000000000000100001010001;
		16'b1111101011000111 : data_out =  24'b000000000000100001010011;
		16'b1111101011001001 : data_out =  24'b000000000000100001010110;
		16'b1111101011001011 : data_out =  24'b000000000000100001011000;
		16'b1111101011001101 : data_out =  24'b000000000000100001011010;
		16'b1111101011001111 : data_out =  24'b000000000000100001011100;
		16'b1111101011010001 : data_out =  24'b000000000000100001011110;
		16'b1111101011010011 : data_out =  24'b000000000000100001100000;
		16'b1111101011010101 : data_out =  24'b000000000000100001100010;
		16'b1111101011011000 : data_out =  24'b000000000000100001100101;
		16'b1111101011011010 : data_out =  24'b000000000000100001100111;
		16'b1111101011011100 : data_out =  24'b000000000000100001101001;
		16'b1111101011011110 : data_out =  24'b000000000000100001101011;
		16'b1111101011100000 : data_out =  24'b000000000000100001101101;
		16'b1111101011100010 : data_out =  24'b000000000000100001101111;
		16'b1111101011100100 : data_out =  24'b000000000000100001110001;
		16'b1111101011100110 : data_out =  24'b000000000000100001110100;
		16'b1111101011101000 : data_out =  24'b000000000000100001110110;
		16'b1111101011101010 : data_out =  24'b000000000000100001111000;
		16'b1111101011101100 : data_out =  24'b000000000000100001111010;
		16'b1111101011101110 : data_out =  24'b000000000000100001111100;
		16'b1111101011110000 : data_out =  24'b000000000000100001111110;
		16'b1111101011110010 : data_out =  24'b000000000000100010000001;
		16'b1111101011110100 : data_out =  24'b000000000000100010000011;
		16'b1111101011110110 : data_out =  24'b000000000000100010000101;
		16'b1111101011111000 : data_out =  24'b000000000000100010000111;
		16'b1111101011111010 : data_out =  24'b000000000000100010001001;
		16'b1111101011111100 : data_out =  24'b000000000000100010001100;
		16'b1111101011111110 : data_out =  24'b000000000000100010001110;
		16'b1111101100000001 : data_out =  24'b000000000000100010010000;
		16'b1111101100000011 : data_out =  24'b000000000000100010010010;
		16'b1111101100000101 : data_out =  24'b000000000000100010010100;
		16'b1111101100000111 : data_out =  24'b000000000000100010010111;
		16'b1111101100001001 : data_out =  24'b000000000000100010011001;
		16'b1111101100001011 : data_out =  24'b000000000000100010011011;
		16'b1111101100001101 : data_out =  24'b000000000000100010011101;
		16'b1111101100001111 : data_out =  24'b000000000000100010011111;
		16'b1111101100010001 : data_out =  24'b000000000000100010100010;
		16'b1111101100010011 : data_out =  24'b000000000000100010100100;
		16'b1111101100010101 : data_out =  24'b000000000000100010100110;
		16'b1111101100010111 : data_out =  24'b000000000000100010101000;
		16'b1111101100011001 : data_out =  24'b000000000000100010101010;
		16'b1111101100011011 : data_out =  24'b000000000000100010101101;
		16'b1111101100011101 : data_out =  24'b000000000000100010101111;
		16'b1111101100011111 : data_out =  24'b000000000000100010110001;
		16'b1111101100100001 : data_out =  24'b000000000000100010110011;
		16'b1111101100100011 : data_out =  24'b000000000000100010110110;
		16'b1111101100100101 : data_out =  24'b000000000000100010111000;
		16'b1111101100100111 : data_out =  24'b000000000000100010111010;
		16'b1111101100101001 : data_out =  24'b000000000000100010111100;
		16'b1111101100101100 : data_out =  24'b000000000000100010111110;
		16'b1111101100101110 : data_out =  24'b000000000000100011000001;
		16'b1111101100110000 : data_out =  24'b000000000000100011000011;
		16'b1111101100110010 : data_out =  24'b000000000000100011000101;
		16'b1111101100110100 : data_out =  24'b000000000000100011000111;
		16'b1111101100110110 : data_out =  24'b000000000000100011001010;
		16'b1111101100111000 : data_out =  24'b000000000000100011001100;
		16'b1111101100111010 : data_out =  24'b000000000000100011001110;
		16'b1111101100111100 : data_out =  24'b000000000000100011010000;
		16'b1111101100111110 : data_out =  24'b000000000000100011010011;
		16'b1111101101000000 : data_out =  24'b000000000000100011010101;
		16'b1111101101000010 : data_out =  24'b000000000000100011010111;
		16'b1111101101000100 : data_out =  24'b000000000000100011011001;
		16'b1111101101000110 : data_out =  24'b000000000000100011011100;
		16'b1111101101001000 : data_out =  24'b000000000000100011011110;
		16'b1111101101001010 : data_out =  24'b000000000000100011100000;
		16'b1111101101001100 : data_out =  24'b000000000000100011100011;
		16'b1111101101001110 : data_out =  24'b000000000000100011100101;
		16'b1111101101010000 : data_out =  24'b000000000000100011100111;
		16'b1111101101010010 : data_out =  24'b000000000000100011101001;
		16'b1111101101010100 : data_out =  24'b000000000000100011101100;
		16'b1111101101010111 : data_out =  24'b000000000000100011101110;
		16'b1111101101011001 : data_out =  24'b000000000000100011110000;
		16'b1111101101011011 : data_out =  24'b000000000000100011110011;
		16'b1111101101011101 : data_out =  24'b000000000000100011110101;
		16'b1111101101011111 : data_out =  24'b000000000000100011110111;
		16'b1111101101100001 : data_out =  24'b000000000000100011111001;
		16'b1111101101100011 : data_out =  24'b000000000000100011111100;
		16'b1111101101100101 : data_out =  24'b000000000000100011111110;
		16'b1111101101100111 : data_out =  24'b000000000000100100000000;
		16'b1111101101101001 : data_out =  24'b000000000000100100000011;
		16'b1111101101101011 : data_out =  24'b000000000000100100000101;
		16'b1111101101101101 : data_out =  24'b000000000000100100000111;
		16'b1111101101101111 : data_out =  24'b000000000000100100001010;
		16'b1111101101110001 : data_out =  24'b000000000000100100001100;
		16'b1111101101110011 : data_out =  24'b000000000000100100001110;
		16'b1111101101110101 : data_out =  24'b000000000000100100010001;
		16'b1111101101110111 : data_out =  24'b000000000000100100010011;
		16'b1111101101111001 : data_out =  24'b000000000000100100010101;
		16'b1111101101111011 : data_out =  24'b000000000000100100011000;
		16'b1111101101111101 : data_out =  24'b000000000000100100011010;
		16'b1111101101111111 : data_out =  24'b000000000000100100011100;
		16'b1111101110000010 : data_out =  24'b000000000000100100011110;
		16'b1111101110000100 : data_out =  24'b000000000000100100100001;
		16'b1111101110000110 : data_out =  24'b000000000000100100100011;
		16'b1111101110001000 : data_out =  24'b000000000000100100100110;
		16'b1111101110001010 : data_out =  24'b000000000000100100101000;
		16'b1111101110001100 : data_out =  24'b000000000000100100101010;
		16'b1111101110001110 : data_out =  24'b000000000000100100101101;
		16'b1111101110010000 : data_out =  24'b000000000000100100101111;
		16'b1111101110010010 : data_out =  24'b000000000000100100110001;
		16'b1111101110010100 : data_out =  24'b000000000000100100110100;
		16'b1111101110010110 : data_out =  24'b000000000000100100110110;
		16'b1111101110011000 : data_out =  24'b000000000000100100111000;
		16'b1111101110011010 : data_out =  24'b000000000000100100111011;
		16'b1111101110011100 : data_out =  24'b000000000000100100111101;
		16'b1111101110011110 : data_out =  24'b000000000000100100111111;
		16'b1111101110100000 : data_out =  24'b000000000000100101000010;
		16'b1111101110100010 : data_out =  24'b000000000000100101000100;
		16'b1111101110100100 : data_out =  24'b000000000000100101000111;
		16'b1111101110100110 : data_out =  24'b000000000000100101001001;
		16'b1111101110101000 : data_out =  24'b000000000000100101001011;
		16'b1111101110101010 : data_out =  24'b000000000000100101001110;
		16'b1111101110101101 : data_out =  24'b000000000000100101010000;
		16'b1111101110101111 : data_out =  24'b000000000000100101010010;
		16'b1111101110110001 : data_out =  24'b000000000000100101010101;
		16'b1111101110110011 : data_out =  24'b000000000000100101010111;
		16'b1111101110110101 : data_out =  24'b000000000000100101011010;
		16'b1111101110110111 : data_out =  24'b000000000000100101011100;
		16'b1111101110111001 : data_out =  24'b000000000000100101011110;
		16'b1111101110111011 : data_out =  24'b000000000000100101100001;
		16'b1111101110111101 : data_out =  24'b000000000000100101100011;
		16'b1111101110111111 : data_out =  24'b000000000000100101100110;
		16'b1111101111000001 : data_out =  24'b000000000000100101101000;
		16'b1111101111000011 : data_out =  24'b000000000000100101101010;
		16'b1111101111000101 : data_out =  24'b000000000000100101101101;
		16'b1111101111000111 : data_out =  24'b000000000000100101101111;
		16'b1111101111001001 : data_out =  24'b000000000000100101110010;
		16'b1111101111001011 : data_out =  24'b000000000000100101110100;
		16'b1111101111001101 : data_out =  24'b000000000000100101110111;
		16'b1111101111001111 : data_out =  24'b000000000000100101111001;
		16'b1111101111010001 : data_out =  24'b000000000000100101111011;
		16'b1111101111010011 : data_out =  24'b000000000000100101111110;
		16'b1111101111010101 : data_out =  24'b000000000000100110000000;
		16'b1111101111011000 : data_out =  24'b000000000000100110000011;
		16'b1111101111011010 : data_out =  24'b000000000000100110000101;
		16'b1111101111011100 : data_out =  24'b000000000000100110001000;
		16'b1111101111011110 : data_out =  24'b000000000000100110001010;
		16'b1111101111100000 : data_out =  24'b000000000000100110001100;
		16'b1111101111100010 : data_out =  24'b000000000000100110001111;
		16'b1111101111100100 : data_out =  24'b000000000000100110010001;
		16'b1111101111100110 : data_out =  24'b000000000000100110010100;
		16'b1111101111101000 : data_out =  24'b000000000000100110010110;
		16'b1111101111101010 : data_out =  24'b000000000000100110011001;
		16'b1111101111101100 : data_out =  24'b000000000000100110011011;
		16'b1111101111101110 : data_out =  24'b000000000000100110011110;
		16'b1111101111110000 : data_out =  24'b000000000000100110100000;
		16'b1111101111110010 : data_out =  24'b000000000000100110100011;
		16'b1111101111110100 : data_out =  24'b000000000000100110100101;
		16'b1111101111110110 : data_out =  24'b000000000000100110100111;
		16'b1111101111111000 : data_out =  24'b000000000000100110101010;
		16'b1111101111111010 : data_out =  24'b000000000000100110101100;
		16'b1111101111111100 : data_out =  24'b000000000000100110101111;
		16'b1111101111111110 : data_out =  24'b000000000000100110110001;
		16'b1111110000000001 : data_out =  24'b000000000000100110110100;
		16'b1111110000000011 : data_out =  24'b000000000000100110110110;
		16'b1111110000000101 : data_out =  24'b000000000000100110111001;
		16'b1111110000000111 : data_out =  24'b000000000000100110111011;
		16'b1111110000001001 : data_out =  24'b000000000000100110111110;
		16'b1111110000001011 : data_out =  24'b000000000000100111000000;
		16'b1111110000001101 : data_out =  24'b000000000000100111000011;
		16'b1111110000001111 : data_out =  24'b000000000000100111000101;
		16'b1111110000010001 : data_out =  24'b000000000000100111001000;
		16'b1111110000010011 : data_out =  24'b000000000000100111001010;
		16'b1111110000010101 : data_out =  24'b000000000000100111001101;
		16'b1111110000010111 : data_out =  24'b000000000000100111001111;
		16'b1111110000011001 : data_out =  24'b000000000000100111010010;
		16'b1111110000011011 : data_out =  24'b000000000000100111010100;
		16'b1111110000011101 : data_out =  24'b000000000000100111010111;
		16'b1111110000011111 : data_out =  24'b000000000000100111011001;
		16'b1111110000100001 : data_out =  24'b000000000000100111011100;
		16'b1111110000100011 : data_out =  24'b000000000000100111011110;
		16'b1111110000100101 : data_out =  24'b000000000000100111100001;
		16'b1111110000100111 : data_out =  24'b000000000000100111100100;
		16'b1111110000101001 : data_out =  24'b000000000000100111100110;
		16'b1111110000101100 : data_out =  24'b000000000000100111101001;
		16'b1111110000101110 : data_out =  24'b000000000000100111101011;
		16'b1111110000110000 : data_out =  24'b000000000000100111101110;
		16'b1111110000110010 : data_out =  24'b000000000000100111110000;
		16'b1111110000110100 : data_out =  24'b000000000000100111110011;
		16'b1111110000110110 : data_out =  24'b000000000000100111110101;
		16'b1111110000111000 : data_out =  24'b000000000000100111111000;
		16'b1111110000111010 : data_out =  24'b000000000000100111111010;
		16'b1111110000111100 : data_out =  24'b000000000000100111111101;
		16'b1111110000111110 : data_out =  24'b000000000000101000000000;
		16'b1111110001000000 : data_out =  24'b000000000000101000000010;
		16'b1111110001000010 : data_out =  24'b000000000000101000000101;
		16'b1111110001000100 : data_out =  24'b000000000000101000000111;
		16'b1111110001000110 : data_out =  24'b000000000000101000001010;
		16'b1111110001001000 : data_out =  24'b000000000000101000001100;
		16'b1111110001001010 : data_out =  24'b000000000000101000001111;
		16'b1111110001001100 : data_out =  24'b000000000000101000010001;
		16'b1111110001001110 : data_out =  24'b000000000000101000010100;
		16'b1111110001010000 : data_out =  24'b000000000000101000010111;
		16'b1111110001010010 : data_out =  24'b000000000000101000011001;
		16'b1111110001010100 : data_out =  24'b000000000000101000011100;
		16'b1111110001010111 : data_out =  24'b000000000000101000011110;
		16'b1111110001011001 : data_out =  24'b000000000000101000100001;
		16'b1111110001011011 : data_out =  24'b000000000000101000100100;
		16'b1111110001011101 : data_out =  24'b000000000000101000100110;
		16'b1111110001011111 : data_out =  24'b000000000000101000101001;
		16'b1111110001100001 : data_out =  24'b000000000000101000101011;
		16'b1111110001100011 : data_out =  24'b000000000000101000101110;
		16'b1111110001100101 : data_out =  24'b000000000000101000110001;
		16'b1111110001100111 : data_out =  24'b000000000000101000110011;
		16'b1111110001101001 : data_out =  24'b000000000000101000110110;
		16'b1111110001101011 : data_out =  24'b000000000000101000111000;
		16'b1111110001101101 : data_out =  24'b000000000000101000111011;
		16'b1111110001101111 : data_out =  24'b000000000000101000111110;
		16'b1111110001110001 : data_out =  24'b000000000000101001000000;
		16'b1111110001110011 : data_out =  24'b000000000000101001000011;
		16'b1111110001110101 : data_out =  24'b000000000000101001000110;
		16'b1111110001110111 : data_out =  24'b000000000000101001001000;
		16'b1111110001111001 : data_out =  24'b000000000000101001001011;
		16'b1111110001111011 : data_out =  24'b000000000000101001001101;
		16'b1111110001111101 : data_out =  24'b000000000000101001010000;
		16'b1111110001111111 : data_out =  24'b000000000000101001010011;
		16'b1111110010000010 : data_out =  24'b000000000000101001010101;
		16'b1111110010000100 : data_out =  24'b000000000000101001011000;
		16'b1111110010000110 : data_out =  24'b000000000000101001011011;
		16'b1111110010001000 : data_out =  24'b000000000000101001011101;
		16'b1111110010001010 : data_out =  24'b000000000000101001100000;
		16'b1111110010001100 : data_out =  24'b000000000000101001100011;
		16'b1111110010001110 : data_out =  24'b000000000000101001100101;
		16'b1111110010010000 : data_out =  24'b000000000000101001101000;
		16'b1111110010010010 : data_out =  24'b000000000000101001101011;
		16'b1111110010010100 : data_out =  24'b000000000000101001101101;
		16'b1111110010010110 : data_out =  24'b000000000000101001110000;
		16'b1111110010011000 : data_out =  24'b000000000000101001110011;
		16'b1111110010011010 : data_out =  24'b000000000000101001110101;
		16'b1111110010011100 : data_out =  24'b000000000000101001111000;
		16'b1111110010011110 : data_out =  24'b000000000000101001111011;
		16'b1111110010100000 : data_out =  24'b000000000000101001111101;
		16'b1111110010100010 : data_out =  24'b000000000000101010000000;
		16'b1111110010100100 : data_out =  24'b000000000000101010000011;
		16'b1111110010100110 : data_out =  24'b000000000000101010000101;
		16'b1111110010101000 : data_out =  24'b000000000000101010001000;
		16'b1111110010101010 : data_out =  24'b000000000000101010001011;
		16'b1111110010101101 : data_out =  24'b000000000000101010001110;
		16'b1111110010101111 : data_out =  24'b000000000000101010010000;
		16'b1111110010110001 : data_out =  24'b000000000000101010010011;
		16'b1111110010110011 : data_out =  24'b000000000000101010010110;
		16'b1111110010110101 : data_out =  24'b000000000000101010011000;
		16'b1111110010110111 : data_out =  24'b000000000000101010011011;
		16'b1111110010111001 : data_out =  24'b000000000000101010011110;
		16'b1111110010111011 : data_out =  24'b000000000000101010100001;
		16'b1111110010111101 : data_out =  24'b000000000000101010100011;
		16'b1111110010111111 : data_out =  24'b000000000000101010100110;
		16'b1111110011000001 : data_out =  24'b000000000000101010101001;
		16'b1111110011000011 : data_out =  24'b000000000000101010101011;
		16'b1111110011000101 : data_out =  24'b000000000000101010101110;
		16'b1111110011000111 : data_out =  24'b000000000000101010110001;
		16'b1111110011001001 : data_out =  24'b000000000000101010110100;
		16'b1111110011001011 : data_out =  24'b000000000000101010110110;
		16'b1111110011001101 : data_out =  24'b000000000000101010111001;
		16'b1111110011001111 : data_out =  24'b000000000000101010111100;
		16'b1111110011010001 : data_out =  24'b000000000000101010111111;
		16'b1111110011010011 : data_out =  24'b000000000000101011000001;
		16'b1111110011010101 : data_out =  24'b000000000000101011000100;
		16'b1111110011011000 : data_out =  24'b000000000000101011000111;
		16'b1111110011011010 : data_out =  24'b000000000000101011001010;
		16'b1111110011011100 : data_out =  24'b000000000000101011001100;
		16'b1111110011011110 : data_out =  24'b000000000000101011001111;
		16'b1111110011100000 : data_out =  24'b000000000000101011010010;
		16'b1111110011100010 : data_out =  24'b000000000000101011010101;
		16'b1111110011100100 : data_out =  24'b000000000000101011010111;
		16'b1111110011100110 : data_out =  24'b000000000000101011011010;
		16'b1111110011101000 : data_out =  24'b000000000000101011011101;
		16'b1111110011101010 : data_out =  24'b000000000000101011100000;
		16'b1111110011101100 : data_out =  24'b000000000000101011100011;
		16'b1111110011101110 : data_out =  24'b000000000000101011100101;
		16'b1111110011110000 : data_out =  24'b000000000000101011101000;
		16'b1111110011110010 : data_out =  24'b000000000000101011101011;
		16'b1111110011110100 : data_out =  24'b000000000000101011101110;
		16'b1111110011110110 : data_out =  24'b000000000000101011110001;
		16'b1111110011111000 : data_out =  24'b000000000000101011110011;
		16'b1111110011111010 : data_out =  24'b000000000000101011110110;
		16'b1111110011111100 : data_out =  24'b000000000000101011111001;
		16'b1111110011111110 : data_out =  24'b000000000000101011111100;
		16'b1111110100000001 : data_out =  24'b000000000000101011111111;
		16'b1111110100000011 : data_out =  24'b000000000000101100000001;
		16'b1111110100000101 : data_out =  24'b000000000000101100000100;
		16'b1111110100000111 : data_out =  24'b000000000000101100000111;
		16'b1111110100001001 : data_out =  24'b000000000000101100001010;
		16'b1111110100001011 : data_out =  24'b000000000000101100001101;
		16'b1111110100001101 : data_out =  24'b000000000000101100010000;
		16'b1111110100001111 : data_out =  24'b000000000000101100010010;
		16'b1111110100010001 : data_out =  24'b000000000000101100010101;
		16'b1111110100010011 : data_out =  24'b000000000000101100011000;
		16'b1111110100010101 : data_out =  24'b000000000000101100011011;
		16'b1111110100010111 : data_out =  24'b000000000000101100011110;
		16'b1111110100011001 : data_out =  24'b000000000000101100100001;
		16'b1111110100011011 : data_out =  24'b000000000000101100100011;
		16'b1111110100011101 : data_out =  24'b000000000000101100100110;
		16'b1111110100011111 : data_out =  24'b000000000000101100101001;
		16'b1111110100100001 : data_out =  24'b000000000000101100101100;
		16'b1111110100100011 : data_out =  24'b000000000000101100101111;
		16'b1111110100100101 : data_out =  24'b000000000000101100110010;
		16'b1111110100100111 : data_out =  24'b000000000000101100110101;
		16'b1111110100101001 : data_out =  24'b000000000000101100111000;
		16'b1111110100101100 : data_out =  24'b000000000000101100111010;
		16'b1111110100101110 : data_out =  24'b000000000000101100111101;
		16'b1111110100110000 : data_out =  24'b000000000000101101000000;
		16'b1111110100110010 : data_out =  24'b000000000000101101000011;
		16'b1111110100110100 : data_out =  24'b000000000000101101000110;
		16'b1111110100110110 : data_out =  24'b000000000000101101001001;
		16'b1111110100111000 : data_out =  24'b000000000000101101001100;
		16'b1111110100111010 : data_out =  24'b000000000000101101001111;
		16'b1111110100111100 : data_out =  24'b000000000000101101010001;
		16'b1111110100111110 : data_out =  24'b000000000000101101010100;
		16'b1111110101000000 : data_out =  24'b000000000000101101010111;
		16'b1111110101000010 : data_out =  24'b000000000000101101011010;
		16'b1111110101000100 : data_out =  24'b000000000000101101011101;
		16'b1111110101000110 : data_out =  24'b000000000000101101100000;
		16'b1111110101001000 : data_out =  24'b000000000000101101100011;
		16'b1111110101001010 : data_out =  24'b000000000000101101100110;
		16'b1111110101001100 : data_out =  24'b000000000000101101101001;
		16'b1111110101001110 : data_out =  24'b000000000000101101101100;
		16'b1111110101010000 : data_out =  24'b000000000000101101101111;
		16'b1111110101010010 : data_out =  24'b000000000000101101110010;
		16'b1111110101010100 : data_out =  24'b000000000000101101110100;
		16'b1111110101010111 : data_out =  24'b000000000000101101110111;
		16'b1111110101011001 : data_out =  24'b000000000000101101111010;
		16'b1111110101011011 : data_out =  24'b000000000000101101111101;
		16'b1111110101011101 : data_out =  24'b000000000000101110000000;
		16'b1111110101011111 : data_out =  24'b000000000000101110000011;
		16'b1111110101100001 : data_out =  24'b000000000000101110000110;
		16'b1111110101100011 : data_out =  24'b000000000000101110001001;
		16'b1111110101100101 : data_out =  24'b000000000000101110001100;
		16'b1111110101100111 : data_out =  24'b000000000000101110001111;
		16'b1111110101101001 : data_out =  24'b000000000000101110010010;
		16'b1111110101101011 : data_out =  24'b000000000000101110010101;
		16'b1111110101101101 : data_out =  24'b000000000000101110011000;
		16'b1111110101101111 : data_out =  24'b000000000000101110011011;
		16'b1111110101110001 : data_out =  24'b000000000000101110011110;
		16'b1111110101110011 : data_out =  24'b000000000000101110100001;
		16'b1111110101110101 : data_out =  24'b000000000000101110100100;
		16'b1111110101110111 : data_out =  24'b000000000000101110100111;
		16'b1111110101111001 : data_out =  24'b000000000000101110101010;
		16'b1111110101111011 : data_out =  24'b000000000000101110101101;
		16'b1111110101111101 : data_out =  24'b000000000000101110110000;
		16'b1111110101111111 : data_out =  24'b000000000000101110110011;
		16'b1111110110000010 : data_out =  24'b000000000000101110110110;
		16'b1111110110000100 : data_out =  24'b000000000000101110111001;
		16'b1111110110000110 : data_out =  24'b000000000000101110111100;
		16'b1111110110001000 : data_out =  24'b000000000000101110111111;
		16'b1111110110001010 : data_out =  24'b000000000000101111000010;
		16'b1111110110001100 : data_out =  24'b000000000000101111000101;
		16'b1111110110001110 : data_out =  24'b000000000000101111001000;
		16'b1111110110010000 : data_out =  24'b000000000000101111001011;
		16'b1111110110010010 : data_out =  24'b000000000000101111001110;
		16'b1111110110010100 : data_out =  24'b000000000000101111010001;
		16'b1111110110010110 : data_out =  24'b000000000000101111010100;
		16'b1111110110011000 : data_out =  24'b000000000000101111010111;
		16'b1111110110011010 : data_out =  24'b000000000000101111011010;
		16'b1111110110011100 : data_out =  24'b000000000000101111011101;
		16'b1111110110011110 : data_out =  24'b000000000000101111100000;
		16'b1111110110100000 : data_out =  24'b000000000000101111100011;
		16'b1111110110100010 : data_out =  24'b000000000000101111100110;
		16'b1111110110100100 : data_out =  24'b000000000000101111101001;
		16'b1111110110100110 : data_out =  24'b000000000000101111101100;
		16'b1111110110101000 : data_out =  24'b000000000000101111101111;
		16'b1111110110101010 : data_out =  24'b000000000000101111110010;
		16'b1111110110101101 : data_out =  24'b000000000000101111110101;
		16'b1111110110101111 : data_out =  24'b000000000000101111111000;
		16'b1111110110110001 : data_out =  24'b000000000000101111111011;
		16'b1111110110110011 : data_out =  24'b000000000000101111111111;
		16'b1111110110110101 : data_out =  24'b000000000000110000000010;
		16'b1111110110110111 : data_out =  24'b000000000000110000000101;
		16'b1111110110111001 : data_out =  24'b000000000000110000001000;
		16'b1111110110111011 : data_out =  24'b000000000000110000001011;
		16'b1111110110111101 : data_out =  24'b000000000000110000001110;
		16'b1111110110111111 : data_out =  24'b000000000000110000010001;
		16'b1111110111000001 : data_out =  24'b000000000000110000010100;
		16'b1111110111000011 : data_out =  24'b000000000000110000010111;
		16'b1111110111000101 : data_out =  24'b000000000000110000011010;
		16'b1111110111000111 : data_out =  24'b000000000000110000011101;
		16'b1111110111001001 : data_out =  24'b000000000000110000100000;
		16'b1111110111001011 : data_out =  24'b000000000000110000100100;
		16'b1111110111001101 : data_out =  24'b000000000000110000100111;
		16'b1111110111001111 : data_out =  24'b000000000000110000101010;
		16'b1111110111010001 : data_out =  24'b000000000000110000101101;
		16'b1111110111010011 : data_out =  24'b000000000000110000110000;
		16'b1111110111010101 : data_out =  24'b000000000000110000110011;
		16'b1111110111011000 : data_out =  24'b000000000000110000110110;
		16'b1111110111011010 : data_out =  24'b000000000000110000111001;
		16'b1111110111011100 : data_out =  24'b000000000000110000111101;
		16'b1111110111011110 : data_out =  24'b000000000000110001000000;
		16'b1111110111100000 : data_out =  24'b000000000000110001000011;
		16'b1111110111100010 : data_out =  24'b000000000000110001000110;
		16'b1111110111100100 : data_out =  24'b000000000000110001001001;
		16'b1111110111100110 : data_out =  24'b000000000000110001001100;
		16'b1111110111101000 : data_out =  24'b000000000000110001001111;
		16'b1111110111101010 : data_out =  24'b000000000000110001010011;
		16'b1111110111101100 : data_out =  24'b000000000000110001010110;
		16'b1111110111101110 : data_out =  24'b000000000000110001011001;
		16'b1111110111110000 : data_out =  24'b000000000000110001011100;
		16'b1111110111110010 : data_out =  24'b000000000000110001011111;
		16'b1111110111110100 : data_out =  24'b000000000000110001100010;
		16'b1111110111110110 : data_out =  24'b000000000000110001100110;
		16'b1111110111111000 : data_out =  24'b000000000000110001101001;
		16'b1111110111111010 : data_out =  24'b000000000000110001101100;
		16'b1111110111111100 : data_out =  24'b000000000000110001101111;
		16'b1111110111111110 : data_out =  24'b000000000000110001110010;
		16'b1111111000000001 : data_out =  24'b000000000000110001110101;
		16'b1111111000000011 : data_out =  24'b000000000000110001111001;
		16'b1111111000000101 : data_out =  24'b000000000000110001111100;
		16'b1111111000000111 : data_out =  24'b000000000000110001111111;
		16'b1111111000001001 : data_out =  24'b000000000000110010000010;
		16'b1111111000001011 : data_out =  24'b000000000000110010000101;
		16'b1111111000001101 : data_out =  24'b000000000000110010001001;
		16'b1111111000001111 : data_out =  24'b000000000000110010001100;
		16'b1111111000010001 : data_out =  24'b000000000000110010001111;
		16'b1111111000010011 : data_out =  24'b000000000000110010010010;
		16'b1111111000010101 : data_out =  24'b000000000000110010010110;
		16'b1111111000010111 : data_out =  24'b000000000000110010011001;
		16'b1111111000011001 : data_out =  24'b000000000000110010011100;
		16'b1111111000011011 : data_out =  24'b000000000000110010011111;
		16'b1111111000011101 : data_out =  24'b000000000000110010100010;
		16'b1111111000011111 : data_out =  24'b000000000000110010100110;
		16'b1111111000100001 : data_out =  24'b000000000000110010101001;
		16'b1111111000100011 : data_out =  24'b000000000000110010101100;
		16'b1111111000100101 : data_out =  24'b000000000000110010101111;
		16'b1111111000100111 : data_out =  24'b000000000000110010110011;
		16'b1111111000101001 : data_out =  24'b000000000000110010110110;
		16'b1111111000101100 : data_out =  24'b000000000000110010111001;
		16'b1111111000101110 : data_out =  24'b000000000000110010111100;
		16'b1111111000110000 : data_out =  24'b000000000000110011000000;
		16'b1111111000110010 : data_out =  24'b000000000000110011000011;
		16'b1111111000110100 : data_out =  24'b000000000000110011000110;
		16'b1111111000110110 : data_out =  24'b000000000000110011001001;
		16'b1111111000111000 : data_out =  24'b000000000000110011001101;
		16'b1111111000111010 : data_out =  24'b000000000000110011010000;
		16'b1111111000111100 : data_out =  24'b000000000000110011010011;
		16'b1111111000111110 : data_out =  24'b000000000000110011010111;
		16'b1111111001000000 : data_out =  24'b000000000000110011011010;
		16'b1111111001000010 : data_out =  24'b000000000000110011011101;
		16'b1111111001000100 : data_out =  24'b000000000000110011100000;
		16'b1111111001000110 : data_out =  24'b000000000000110011100100;
		16'b1111111001001000 : data_out =  24'b000000000000110011100111;
		16'b1111111001001010 : data_out =  24'b000000000000110011101010;
		16'b1111111001001100 : data_out =  24'b000000000000110011101110;
		16'b1111111001001110 : data_out =  24'b000000000000110011110001;
		16'b1111111001010000 : data_out =  24'b000000000000110011110100;
		16'b1111111001010010 : data_out =  24'b000000000000110011111000;
		16'b1111111001010100 : data_out =  24'b000000000000110011111011;
		16'b1111111001010111 : data_out =  24'b000000000000110011111110;
		16'b1111111001011001 : data_out =  24'b000000000000110100000010;
		16'b1111111001011011 : data_out =  24'b000000000000110100000101;
		16'b1111111001011101 : data_out =  24'b000000000000110100001000;
		16'b1111111001011111 : data_out =  24'b000000000000110100001100;
		16'b1111111001100001 : data_out =  24'b000000000000110100001111;
		16'b1111111001100011 : data_out =  24'b000000000000110100010010;
		16'b1111111001100101 : data_out =  24'b000000000000110100010110;
		16'b1111111001100111 : data_out =  24'b000000000000110100011001;
		16'b1111111001101001 : data_out =  24'b000000000000110100011100;
		16'b1111111001101011 : data_out =  24'b000000000000110100100000;
		16'b1111111001101101 : data_out =  24'b000000000000110100100011;
		16'b1111111001101111 : data_out =  24'b000000000000110100100110;
		16'b1111111001110001 : data_out =  24'b000000000000110100101010;
		16'b1111111001110011 : data_out =  24'b000000000000110100101101;
		16'b1111111001110101 : data_out =  24'b000000000000110100110001;
		16'b1111111001110111 : data_out =  24'b000000000000110100110100;
		16'b1111111001111001 : data_out =  24'b000000000000110100110111;
		16'b1111111001111011 : data_out =  24'b000000000000110100111011;
		16'b1111111001111101 : data_out =  24'b000000000000110100111110;
		16'b1111111001111111 : data_out =  24'b000000000000110101000010;
		16'b1111111010000010 : data_out =  24'b000000000000110101000101;
		16'b1111111010000100 : data_out =  24'b000000000000110101001000;
		16'b1111111010000110 : data_out =  24'b000000000000110101001100;
		16'b1111111010001000 : data_out =  24'b000000000000110101001111;
		16'b1111111010001010 : data_out =  24'b000000000000110101010011;
		16'b1111111010001100 : data_out =  24'b000000000000110101010110;
		16'b1111111010001110 : data_out =  24'b000000000000110101011001;
		16'b1111111010010000 : data_out =  24'b000000000000110101011101;
		16'b1111111010010010 : data_out =  24'b000000000000110101100000;
		16'b1111111010010100 : data_out =  24'b000000000000110101100100;
		16'b1111111010010110 : data_out =  24'b000000000000110101100111;
		16'b1111111010011000 : data_out =  24'b000000000000110101101010;
		16'b1111111010011010 : data_out =  24'b000000000000110101101110;
		16'b1111111010011100 : data_out =  24'b000000000000110101110001;
		16'b1111111010011110 : data_out =  24'b000000000000110101110101;
		16'b1111111010100000 : data_out =  24'b000000000000110101111000;
		16'b1111111010100010 : data_out =  24'b000000000000110101111100;
		16'b1111111010100100 : data_out =  24'b000000000000110101111111;
		16'b1111111010100110 : data_out =  24'b000000000000110110000011;
		16'b1111111010101000 : data_out =  24'b000000000000110110000110;
		16'b1111111010101010 : data_out =  24'b000000000000110110001010;
		16'b1111111010101101 : data_out =  24'b000000000000110110001101;
		16'b1111111010101111 : data_out =  24'b000000000000110110010000;
		16'b1111111010110001 : data_out =  24'b000000000000110110010100;
		16'b1111111010110011 : data_out =  24'b000000000000110110010111;
		16'b1111111010110101 : data_out =  24'b000000000000110110011011;
		16'b1111111010110111 : data_out =  24'b000000000000110110011110;
		16'b1111111010111001 : data_out =  24'b000000000000110110100010;
		16'b1111111010111011 : data_out =  24'b000000000000110110100101;
		16'b1111111010111101 : data_out =  24'b000000000000110110101001;
		16'b1111111010111111 : data_out =  24'b000000000000110110101100;
		16'b1111111011000001 : data_out =  24'b000000000000110110110000;
		16'b1111111011000011 : data_out =  24'b000000000000110110110011;
		16'b1111111011000101 : data_out =  24'b000000000000110110110111;
		16'b1111111011000111 : data_out =  24'b000000000000110110111010;
		16'b1111111011001001 : data_out =  24'b000000000000110110111110;
		16'b1111111011001011 : data_out =  24'b000000000000110111000001;
		16'b1111111011001101 : data_out =  24'b000000000000110111000101;
		16'b1111111011001111 : data_out =  24'b000000000000110111001000;
		16'b1111111011010001 : data_out =  24'b000000000000110111001100;
		16'b1111111011010011 : data_out =  24'b000000000000110111010000;
		16'b1111111011010101 : data_out =  24'b000000000000110111010011;
		16'b1111111011011000 : data_out =  24'b000000000000110111010111;
		16'b1111111011011010 : data_out =  24'b000000000000110111011010;
		16'b1111111011011100 : data_out =  24'b000000000000110111011110;
		16'b1111111011011110 : data_out =  24'b000000000000110111100001;
		16'b1111111011100000 : data_out =  24'b000000000000110111100101;
		16'b1111111011100010 : data_out =  24'b000000000000110111101000;
		16'b1111111011100100 : data_out =  24'b000000000000110111101100;
		16'b1111111011100110 : data_out =  24'b000000000000110111110000;
		16'b1111111011101000 : data_out =  24'b000000000000110111110011;
		16'b1111111011101010 : data_out =  24'b000000000000110111110111;
		16'b1111111011101100 : data_out =  24'b000000000000110111111010;
		16'b1111111011101110 : data_out =  24'b000000000000110111111110;
		16'b1111111011110000 : data_out =  24'b000000000000111000000001;
		16'b1111111011110010 : data_out =  24'b000000000000111000000101;
		16'b1111111011110100 : data_out =  24'b000000000000111000001001;
		16'b1111111011110110 : data_out =  24'b000000000000111000001100;
		16'b1111111011111000 : data_out =  24'b000000000000111000010000;
		16'b1111111011111010 : data_out =  24'b000000000000111000010011;
		16'b1111111011111100 : data_out =  24'b000000000000111000010111;
		16'b1111111011111110 : data_out =  24'b000000000000111000011011;
		16'b1111111100000001 : data_out =  24'b000000000000111000011110;
		16'b1111111100000011 : data_out =  24'b000000000000111000100010;
		16'b1111111100000101 : data_out =  24'b000000000000111000100101;
		16'b1111111100000111 : data_out =  24'b000000000000111000101001;
		16'b1111111100001001 : data_out =  24'b000000000000111000101101;
		16'b1111111100001011 : data_out =  24'b000000000000111000110000;
		16'b1111111100001101 : data_out =  24'b000000000000111000110100;
		16'b1111111100001111 : data_out =  24'b000000000000111000111000;
		16'b1111111100010001 : data_out =  24'b000000000000111000111011;
		16'b1111111100010011 : data_out =  24'b000000000000111000111111;
		16'b1111111100010101 : data_out =  24'b000000000000111001000011;
		16'b1111111100010111 : data_out =  24'b000000000000111001000110;
		16'b1111111100011001 : data_out =  24'b000000000000111001001010;
		16'b1111111100011011 : data_out =  24'b000000000000111001001110;
		16'b1111111100011101 : data_out =  24'b000000000000111001010001;
		16'b1111111100011111 : data_out =  24'b000000000000111001010101;
		16'b1111111100100001 : data_out =  24'b000000000000111001011001;
		16'b1111111100100011 : data_out =  24'b000000000000111001011100;
		16'b1111111100100101 : data_out =  24'b000000000000111001100000;
		16'b1111111100100111 : data_out =  24'b000000000000111001100100;
		16'b1111111100101001 : data_out =  24'b000000000000111001100111;
		16'b1111111100101100 : data_out =  24'b000000000000111001101011;
		16'b1111111100101110 : data_out =  24'b000000000000111001101111;
		16'b1111111100110000 : data_out =  24'b000000000000111001110010;
		16'b1111111100110010 : data_out =  24'b000000000000111001110110;
		16'b1111111100110100 : data_out =  24'b000000000000111001111010;
		16'b1111111100110110 : data_out =  24'b000000000000111001111101;
		16'b1111111100111000 : data_out =  24'b000000000000111010000001;
		16'b1111111100111010 : data_out =  24'b000000000000111010000101;
		16'b1111111100111100 : data_out =  24'b000000000000111010001001;
		16'b1111111100111110 : data_out =  24'b000000000000111010001100;
		16'b1111111101000000 : data_out =  24'b000000000000111010010000;
		16'b1111111101000010 : data_out =  24'b000000000000111010010100;
		16'b1111111101000100 : data_out =  24'b000000000000111010010111;
		16'b1111111101000110 : data_out =  24'b000000000000111010011011;
		16'b1111111101001000 : data_out =  24'b000000000000111010011111;
		16'b1111111101001010 : data_out =  24'b000000000000111010100011;
		16'b1111111101001100 : data_out =  24'b000000000000111010100110;
		16'b1111111101001110 : data_out =  24'b000000000000111010101010;
		16'b1111111101010000 : data_out =  24'b000000000000111010101110;
		16'b1111111101010010 : data_out =  24'b000000000000111010110010;
		16'b1111111101010100 : data_out =  24'b000000000000111010110101;
		16'b1111111101010111 : data_out =  24'b000000000000111010111001;
		16'b1111111101011001 : data_out =  24'b000000000000111010111101;
		16'b1111111101011011 : data_out =  24'b000000000000111011000001;
		16'b1111111101011101 : data_out =  24'b000000000000111011000101;
		16'b1111111101011111 : data_out =  24'b000000000000111011001000;
		16'b1111111101100001 : data_out =  24'b000000000000111011001100;
		16'b1111111101100011 : data_out =  24'b000000000000111011010000;
		16'b1111111101100101 : data_out =  24'b000000000000111011010100;
		16'b1111111101100111 : data_out =  24'b000000000000111011011000;
		16'b1111111101101001 : data_out =  24'b000000000000111011011011;
		16'b1111111101101011 : data_out =  24'b000000000000111011011111;
		16'b1111111101101101 : data_out =  24'b000000000000111011100011;
		16'b1111111101101111 : data_out =  24'b000000000000111011100111;
		16'b1111111101110001 : data_out =  24'b000000000000111011101011;
		16'b1111111101110011 : data_out =  24'b000000000000111011101110;
		16'b1111111101110101 : data_out =  24'b000000000000111011110010;
		16'b1111111101110111 : data_out =  24'b000000000000111011110110;
		16'b1111111101111001 : data_out =  24'b000000000000111011111010;
		16'b1111111101111011 : data_out =  24'b000000000000111011111110;
		16'b1111111101111101 : data_out =  24'b000000000000111100000010;
		16'b1111111101111111 : data_out =  24'b000000000000111100000101;
		16'b1111111110000010 : data_out =  24'b000000000000111100001001;
		16'b1111111110000100 : data_out =  24'b000000000000111100001101;
		16'b1111111110000110 : data_out =  24'b000000000000111100010001;
		16'b1111111110001000 : data_out =  24'b000000000000111100010101;
		16'b1111111110001010 : data_out =  24'b000000000000111100011001;
		16'b1111111110001100 : data_out =  24'b000000000000111100011101;
		16'b1111111110001110 : data_out =  24'b000000000000111100100000;
		16'b1111111110010000 : data_out =  24'b000000000000111100100100;
		16'b1111111110010010 : data_out =  24'b000000000000111100101000;
		16'b1111111110010100 : data_out =  24'b000000000000111100101100;
		16'b1111111110010110 : data_out =  24'b000000000000111100110000;
		16'b1111111110011000 : data_out =  24'b000000000000111100110100;
		16'b1111111110011010 : data_out =  24'b000000000000111100111000;
		16'b1111111110011100 : data_out =  24'b000000000000111100111100;
		16'b1111111110011110 : data_out =  24'b000000000000111101000000;
		16'b1111111110100000 : data_out =  24'b000000000000111101000011;
		16'b1111111110100010 : data_out =  24'b000000000000111101000111;
		16'b1111111110100100 : data_out =  24'b000000000000111101001011;
		16'b1111111110100110 : data_out =  24'b000000000000111101001111;
		16'b1111111110101000 : data_out =  24'b000000000000111101010011;
		16'b1111111110101010 : data_out =  24'b000000000000111101010111;
		16'b1111111110101101 : data_out =  24'b000000000000111101011011;
		16'b1111111110101111 : data_out =  24'b000000000000111101011111;
		16'b1111111110110001 : data_out =  24'b000000000000111101100011;
		16'b1111111110110011 : data_out =  24'b000000000000111101100111;
		16'b1111111110110101 : data_out =  24'b000000000000111101101011;
		16'b1111111110110111 : data_out =  24'b000000000000111101101111;
		16'b1111111110111001 : data_out =  24'b000000000000111101110011;
		16'b1111111110111011 : data_out =  24'b000000000000111101110111;
		16'b1111111110111101 : data_out =  24'b000000000000111101111011;
		16'b1111111110111111 : data_out =  24'b000000000000111101111111;
		16'b1111111111000001 : data_out =  24'b000000000000111110000010;
		16'b1111111111000011 : data_out =  24'b000000000000111110000110;
		16'b1111111111000101 : data_out =  24'b000000000000111110001010;
		16'b1111111111000111 : data_out =  24'b000000000000111110001110;
		16'b1111111111001001 : data_out =  24'b000000000000111110010010;
		16'b1111111111001011 : data_out =  24'b000000000000111110010110;
		16'b1111111111001101 : data_out =  24'b000000000000111110011010;
		16'b1111111111001111 : data_out =  24'b000000000000111110011110;
		16'b1111111111010001 : data_out =  24'b000000000000111110100010;
		16'b1111111111010011 : data_out =  24'b000000000000111110100110;
		16'b1111111111010101 : data_out =  24'b000000000000111110101010;
		16'b1111111111011000 : data_out =  24'b000000000000111110101110;
		16'b1111111111011010 : data_out =  24'b000000000000111110110010;
		16'b1111111111011100 : data_out =  24'b000000000000111110110110;
		16'b1111111111011110 : data_out =  24'b000000000000111110111010;
		16'b1111111111100000 : data_out =  24'b000000000000111110111110;
		16'b1111111111100010 : data_out =  24'b000000000000111111000011;
		16'b1111111111100100 : data_out =  24'b000000000000111111000111;
		16'b1111111111100110 : data_out =  24'b000000000000111111001011;
		16'b1111111111101000 : data_out =  24'b000000000000111111001111;
		16'b1111111111101010 : data_out =  24'b000000000000111111010011;
		16'b1111111111101100 : data_out =  24'b000000000000111111010111;
		16'b1111111111101110 : data_out =  24'b000000000000111111011011;
		16'b1111111111110000 : data_out =  24'b000000000000111111011111;
		16'b1111111111110010 : data_out =  24'b000000000000111111100011;
		16'b1111111111110100 : data_out =  24'b000000000000111111100111;
		16'b1111111111110110 : data_out =  24'b000000000000111111101011;
		16'b1111111111111000 : data_out =  24'b000000000000111111101111;
		16'b1111111111111010 : data_out =  24'b000000000000111111110011;
		16'b1111111111111100 : data_out =  24'b000000000000111111110111;
		16'b1111111111111110 : data_out =  24'b000000000000111111111011;
		16'b0000000000000000 : data_out =  24'b000000000001000000000000;
		16'b0000000000000010 : data_out =  24'b000000000001000000000100;
		16'b0000000000000100 : data_out =  24'b000000000001000000001000;
		16'b0000000000000110 : data_out =  24'b000000000001000000001100;
		16'b0000000000001000 : data_out =  24'b000000000001000000010000;
		16'b0000000000001010 : data_out =  24'b000000000001000000010100;
		16'b0000000000001100 : data_out =  24'b000000000001000000011000;
		16'b0000000000001110 : data_out =  24'b000000000001000000011100;
		16'b0000000000010000 : data_out =  24'b000000000001000000100000;
		16'b0000000000010010 : data_out =  24'b000000000001000000100101;
		16'b0000000000010100 : data_out =  24'b000000000001000000101001;
		16'b0000000000010110 : data_out =  24'b000000000001000000101101;
		16'b0000000000011000 : data_out =  24'b000000000001000000110001;
		16'b0000000000011010 : data_out =  24'b000000000001000000110101;
		16'b0000000000011100 : data_out =  24'b000000000001000000111001;
		16'b0000000000011110 : data_out =  24'b000000000001000000111101;
		16'b0000000000100000 : data_out =  24'b000000000001000001000010;
		16'b0000000000100010 : data_out =  24'b000000000001000001000110;
		16'b0000000000100100 : data_out =  24'b000000000001000001001010;
		16'b0000000000100110 : data_out =  24'b000000000001000001001110;
		16'b0000000000101000 : data_out =  24'b000000000001000001010010;
		16'b0000000000101011 : data_out =  24'b000000000001000001010110;
		16'b0000000000101101 : data_out =  24'b000000000001000001011011;
		16'b0000000000101111 : data_out =  24'b000000000001000001011111;
		16'b0000000000110001 : data_out =  24'b000000000001000001100011;
		16'b0000000000110011 : data_out =  24'b000000000001000001100111;
		16'b0000000000110101 : data_out =  24'b000000000001000001101011;
		16'b0000000000110111 : data_out =  24'b000000000001000001110000;
		16'b0000000000111001 : data_out =  24'b000000000001000001110100;
		16'b0000000000111011 : data_out =  24'b000000000001000001111000;
		16'b0000000000111101 : data_out =  24'b000000000001000001111100;
		16'b0000000000111111 : data_out =  24'b000000000001000010000000;
		16'b0000000001000001 : data_out =  24'b000000000001000010000101;
		16'b0000000001000011 : data_out =  24'b000000000001000010001001;
		16'b0000000001000101 : data_out =  24'b000000000001000010001101;
		16'b0000000001000111 : data_out =  24'b000000000001000010010001;
		16'b0000000001001001 : data_out =  24'b000000000001000010010110;
		16'b0000000001001011 : data_out =  24'b000000000001000010011010;
		16'b0000000001001101 : data_out =  24'b000000000001000010011110;
		16'b0000000001001111 : data_out =  24'b000000000001000010100010;
		16'b0000000001010001 : data_out =  24'b000000000001000010100111;
		16'b0000000001010011 : data_out =  24'b000000000001000010101011;
		16'b0000000001010110 : data_out =  24'b000000000001000010101111;
		16'b0000000001011000 : data_out =  24'b000000000001000010110011;
		16'b0000000001011010 : data_out =  24'b000000000001000010111000;
		16'b0000000001011100 : data_out =  24'b000000000001000010111100;
		16'b0000000001011110 : data_out =  24'b000000000001000011000000;
		16'b0000000001100000 : data_out =  24'b000000000001000011000101;
		16'b0000000001100010 : data_out =  24'b000000000001000011001001;
		16'b0000000001100100 : data_out =  24'b000000000001000011001101;
		16'b0000000001100110 : data_out =  24'b000000000001000011010010;
		16'b0000000001101000 : data_out =  24'b000000000001000011010110;
		16'b0000000001101010 : data_out =  24'b000000000001000011011010;
		16'b0000000001101100 : data_out =  24'b000000000001000011011110;
		16'b0000000001101110 : data_out =  24'b000000000001000011100011;
		16'b0000000001110000 : data_out =  24'b000000000001000011100111;
		16'b0000000001110010 : data_out =  24'b000000000001000011101011;
		16'b0000000001110100 : data_out =  24'b000000000001000011110000;
		16'b0000000001110110 : data_out =  24'b000000000001000011110100;
		16'b0000000001111000 : data_out =  24'b000000000001000011111000;
		16'b0000000001111010 : data_out =  24'b000000000001000011111101;
		16'b0000000001111100 : data_out =  24'b000000000001000100000001;
		16'b0000000001111110 : data_out =  24'b000000000001000100000101;
		16'b0000000010000001 : data_out =  24'b000000000001000100001010;
		16'b0000000010000011 : data_out =  24'b000000000001000100001110;
		16'b0000000010000101 : data_out =  24'b000000000001000100010011;
		16'b0000000010000111 : data_out =  24'b000000000001000100010111;
		16'b0000000010001001 : data_out =  24'b000000000001000100011011;
		16'b0000000010001011 : data_out =  24'b000000000001000100100000;
		16'b0000000010001101 : data_out =  24'b000000000001000100100100;
		16'b0000000010001111 : data_out =  24'b000000000001000100101000;
		16'b0000000010010001 : data_out =  24'b000000000001000100101101;
		16'b0000000010010011 : data_out =  24'b000000000001000100110001;
		16'b0000000010010101 : data_out =  24'b000000000001000100110110;
		16'b0000000010010111 : data_out =  24'b000000000001000100111010;
		16'b0000000010011001 : data_out =  24'b000000000001000100111111;
		16'b0000000010011011 : data_out =  24'b000000000001000101000011;
		16'b0000000010011101 : data_out =  24'b000000000001000101000111;
		16'b0000000010011111 : data_out =  24'b000000000001000101001100;
		16'b0000000010100001 : data_out =  24'b000000000001000101010000;
		16'b0000000010100011 : data_out =  24'b000000000001000101010101;
		16'b0000000010100101 : data_out =  24'b000000000001000101011001;
		16'b0000000010100111 : data_out =  24'b000000000001000101011110;
		16'b0000000010101001 : data_out =  24'b000000000001000101100010;
		16'b0000000010101100 : data_out =  24'b000000000001000101100110;
		16'b0000000010101110 : data_out =  24'b000000000001000101101011;
		16'b0000000010110000 : data_out =  24'b000000000001000101101111;
		16'b0000000010110010 : data_out =  24'b000000000001000101110100;
		16'b0000000010110100 : data_out =  24'b000000000001000101111000;
		16'b0000000010110110 : data_out =  24'b000000000001000101111101;
		16'b0000000010111000 : data_out =  24'b000000000001000110000001;
		16'b0000000010111010 : data_out =  24'b000000000001000110000110;
		16'b0000000010111100 : data_out =  24'b000000000001000110001010;
		16'b0000000010111110 : data_out =  24'b000000000001000110001111;
		16'b0000000011000000 : data_out =  24'b000000000001000110010011;
		16'b0000000011000010 : data_out =  24'b000000000001000110011000;
		16'b0000000011000100 : data_out =  24'b000000000001000110011100;
		16'b0000000011000110 : data_out =  24'b000000000001000110100001;
		16'b0000000011001000 : data_out =  24'b000000000001000110100101;
		16'b0000000011001010 : data_out =  24'b000000000001000110101010;
		16'b0000000011001100 : data_out =  24'b000000000001000110101110;
		16'b0000000011001110 : data_out =  24'b000000000001000110110011;
		16'b0000000011010000 : data_out =  24'b000000000001000110110111;
		16'b0000000011010010 : data_out =  24'b000000000001000110111100;
		16'b0000000011010100 : data_out =  24'b000000000001000111000000;
		16'b0000000011010111 : data_out =  24'b000000000001000111000101;
		16'b0000000011011001 : data_out =  24'b000000000001000111001010;
		16'b0000000011011011 : data_out =  24'b000000000001000111001110;
		16'b0000000011011101 : data_out =  24'b000000000001000111010011;
		16'b0000000011011111 : data_out =  24'b000000000001000111010111;
		16'b0000000011100001 : data_out =  24'b000000000001000111011100;
		16'b0000000011100011 : data_out =  24'b000000000001000111100000;
		16'b0000000011100101 : data_out =  24'b000000000001000111100101;
		16'b0000000011100111 : data_out =  24'b000000000001000111101010;
		16'b0000000011101001 : data_out =  24'b000000000001000111101110;
		16'b0000000011101011 : data_out =  24'b000000000001000111110011;
		16'b0000000011101101 : data_out =  24'b000000000001000111110111;
		16'b0000000011101111 : data_out =  24'b000000000001000111111100;
		16'b0000000011110001 : data_out =  24'b000000000001001000000000;
		16'b0000000011110011 : data_out =  24'b000000000001001000000101;
		16'b0000000011110101 : data_out =  24'b000000000001001000001010;
		16'b0000000011110111 : data_out =  24'b000000000001001000001110;
		16'b0000000011111001 : data_out =  24'b000000000001001000010011;
		16'b0000000011111011 : data_out =  24'b000000000001001000011000;
		16'b0000000011111101 : data_out =  24'b000000000001001000011100;
		16'b0000000100000000 : data_out =  24'b000000000001001000100001;
		16'b0000000100000010 : data_out =  24'b000000000001001000100110;
		16'b0000000100000100 : data_out =  24'b000000000001001000101010;
		16'b0000000100000110 : data_out =  24'b000000000001001000101111;
		16'b0000000100001000 : data_out =  24'b000000000001001000110011;
		16'b0000000100001010 : data_out =  24'b000000000001001000111000;
		16'b0000000100001100 : data_out =  24'b000000000001001000111101;
		16'b0000000100001110 : data_out =  24'b000000000001001001000001;
		16'b0000000100010000 : data_out =  24'b000000000001001001000110;
		16'b0000000100010010 : data_out =  24'b000000000001001001001011;
		16'b0000000100010100 : data_out =  24'b000000000001001001010000;
		16'b0000000100010110 : data_out =  24'b000000000001001001010100;
		16'b0000000100011000 : data_out =  24'b000000000001001001011001;
		16'b0000000100011010 : data_out =  24'b000000000001001001011110;
		16'b0000000100011100 : data_out =  24'b000000000001001001100010;
		16'b0000000100011110 : data_out =  24'b000000000001001001100111;
		16'b0000000100100000 : data_out =  24'b000000000001001001101100;
		16'b0000000100100010 : data_out =  24'b000000000001001001110000;
		16'b0000000100100100 : data_out =  24'b000000000001001001110101;
		16'b0000000100100110 : data_out =  24'b000000000001001001111010;
		16'b0000000100101000 : data_out =  24'b000000000001001001111111;
		16'b0000000100101011 : data_out =  24'b000000000001001010000011;
		16'b0000000100101101 : data_out =  24'b000000000001001010001000;
		16'b0000000100101111 : data_out =  24'b000000000001001010001101;
		16'b0000000100110001 : data_out =  24'b000000000001001010010010;
		16'b0000000100110011 : data_out =  24'b000000000001001010010110;
		16'b0000000100110101 : data_out =  24'b000000000001001010011011;
		16'b0000000100110111 : data_out =  24'b000000000001001010100000;
		16'b0000000100111001 : data_out =  24'b000000000001001010100101;
		16'b0000000100111011 : data_out =  24'b000000000001001010101001;
		16'b0000000100111101 : data_out =  24'b000000000001001010101110;
		16'b0000000100111111 : data_out =  24'b000000000001001010110011;
		16'b0000000101000001 : data_out =  24'b000000000001001010111000;
		16'b0000000101000011 : data_out =  24'b000000000001001010111101;
		16'b0000000101000101 : data_out =  24'b000000000001001011000001;
		16'b0000000101000111 : data_out =  24'b000000000001001011000110;
		16'b0000000101001001 : data_out =  24'b000000000001001011001011;
		16'b0000000101001011 : data_out =  24'b000000000001001011010000;
		16'b0000000101001101 : data_out =  24'b000000000001001011010101;
		16'b0000000101001111 : data_out =  24'b000000000001001011011001;
		16'b0000000101010001 : data_out =  24'b000000000001001011011110;
		16'b0000000101010011 : data_out =  24'b000000000001001011100011;
		16'b0000000101010110 : data_out =  24'b000000000001001011101000;
		16'b0000000101011000 : data_out =  24'b000000000001001011101101;
		16'b0000000101011010 : data_out =  24'b000000000001001011110010;
		16'b0000000101011100 : data_out =  24'b000000000001001011110111;
		16'b0000000101011110 : data_out =  24'b000000000001001011111011;
		16'b0000000101100000 : data_out =  24'b000000000001001100000000;
		16'b0000000101100010 : data_out =  24'b000000000001001100000101;
		16'b0000000101100100 : data_out =  24'b000000000001001100001010;
		16'b0000000101100110 : data_out =  24'b000000000001001100001111;
		16'b0000000101101000 : data_out =  24'b000000000001001100010100;
		16'b0000000101101010 : data_out =  24'b000000000001001100011001;
		16'b0000000101101100 : data_out =  24'b000000000001001100011110;
		16'b0000000101101110 : data_out =  24'b000000000001001100100010;
		16'b0000000101110000 : data_out =  24'b000000000001001100100111;
		16'b0000000101110010 : data_out =  24'b000000000001001100101100;
		16'b0000000101110100 : data_out =  24'b000000000001001100110001;
		16'b0000000101110110 : data_out =  24'b000000000001001100110110;
		16'b0000000101111000 : data_out =  24'b000000000001001100111011;
		16'b0000000101111010 : data_out =  24'b000000000001001101000000;
		16'b0000000101111100 : data_out =  24'b000000000001001101000101;
		16'b0000000101111110 : data_out =  24'b000000000001001101001010;
		16'b0000000110000001 : data_out =  24'b000000000001001101001111;
		16'b0000000110000011 : data_out =  24'b000000000001001101010100;
		16'b0000000110000101 : data_out =  24'b000000000001001101011001;
		16'b0000000110000111 : data_out =  24'b000000000001001101011110;
		16'b0000000110001001 : data_out =  24'b000000000001001101100011;
		16'b0000000110001011 : data_out =  24'b000000000001001101100111;
		16'b0000000110001101 : data_out =  24'b000000000001001101101100;
		16'b0000000110001111 : data_out =  24'b000000000001001101110001;
		16'b0000000110010001 : data_out =  24'b000000000001001101110110;
		16'b0000000110010011 : data_out =  24'b000000000001001101111011;
		16'b0000000110010101 : data_out =  24'b000000000001001110000000;
		16'b0000000110010111 : data_out =  24'b000000000001001110000101;
		16'b0000000110011001 : data_out =  24'b000000000001001110001010;
		16'b0000000110011011 : data_out =  24'b000000000001001110001111;
		16'b0000000110011101 : data_out =  24'b000000000001001110010100;
		16'b0000000110011111 : data_out =  24'b000000000001001110011001;
		16'b0000000110100001 : data_out =  24'b000000000001001110011110;
		16'b0000000110100011 : data_out =  24'b000000000001001110100011;
		16'b0000000110100101 : data_out =  24'b000000000001001110101000;
		16'b0000000110100111 : data_out =  24'b000000000001001110101110;
		16'b0000000110101001 : data_out =  24'b000000000001001110110011;
		16'b0000000110101100 : data_out =  24'b000000000001001110111000;
		16'b0000000110101110 : data_out =  24'b000000000001001110111101;
		16'b0000000110110000 : data_out =  24'b000000000001001111000010;
		16'b0000000110110010 : data_out =  24'b000000000001001111000111;
		16'b0000000110110100 : data_out =  24'b000000000001001111001100;
		16'b0000000110110110 : data_out =  24'b000000000001001111010001;
		16'b0000000110111000 : data_out =  24'b000000000001001111010110;
		16'b0000000110111010 : data_out =  24'b000000000001001111011011;
		16'b0000000110111100 : data_out =  24'b000000000001001111100000;
		16'b0000000110111110 : data_out =  24'b000000000001001111100101;
		16'b0000000111000000 : data_out =  24'b000000000001001111101010;
		16'b0000000111000010 : data_out =  24'b000000000001001111101111;
		16'b0000000111000100 : data_out =  24'b000000000001001111110101;
		16'b0000000111000110 : data_out =  24'b000000000001001111111010;
		16'b0000000111001000 : data_out =  24'b000000000001001111111111;
		16'b0000000111001010 : data_out =  24'b000000000001010000000100;
		16'b0000000111001100 : data_out =  24'b000000000001010000001001;
		16'b0000000111001110 : data_out =  24'b000000000001010000001110;
		16'b0000000111010000 : data_out =  24'b000000000001010000010011;
		16'b0000000111010010 : data_out =  24'b000000000001010000011000;
		16'b0000000111010100 : data_out =  24'b000000000001010000011110;
		16'b0000000111010111 : data_out =  24'b000000000001010000100011;
		16'b0000000111011001 : data_out =  24'b000000000001010000101000;
		16'b0000000111011011 : data_out =  24'b000000000001010000101101;
		16'b0000000111011101 : data_out =  24'b000000000001010000110010;
		16'b0000000111011111 : data_out =  24'b000000000001010000110111;
		16'b0000000111100001 : data_out =  24'b000000000001010000111101;
		16'b0000000111100011 : data_out =  24'b000000000001010001000010;
		16'b0000000111100101 : data_out =  24'b000000000001010001000111;
		16'b0000000111100111 : data_out =  24'b000000000001010001001100;
		16'b0000000111101001 : data_out =  24'b000000000001010001010001;
		16'b0000000111101011 : data_out =  24'b000000000001010001010111;
		16'b0000000111101101 : data_out =  24'b000000000001010001011100;
		16'b0000000111101111 : data_out =  24'b000000000001010001100001;
		16'b0000000111110001 : data_out =  24'b000000000001010001100110;
		16'b0000000111110011 : data_out =  24'b000000000001010001101011;
		16'b0000000111110101 : data_out =  24'b000000000001010001110001;
		16'b0000000111110111 : data_out =  24'b000000000001010001110110;
		16'b0000000111111001 : data_out =  24'b000000000001010001111011;
		16'b0000000111111011 : data_out =  24'b000000000001010010000000;
		16'b0000000111111101 : data_out =  24'b000000000001010010000110;
		16'b0000001000000000 : data_out =  24'b000000000001010010001011;
		16'b0000001000000010 : data_out =  24'b000000000001010010010000;
		16'b0000001000000100 : data_out =  24'b000000000001010010010101;
		16'b0000001000000110 : data_out =  24'b000000000001010010011011;
		16'b0000001000001000 : data_out =  24'b000000000001010010100000;
		16'b0000001000001010 : data_out =  24'b000000000001010010100101;
		16'b0000001000001100 : data_out =  24'b000000000001010010101011;
		16'b0000001000001110 : data_out =  24'b000000000001010010110000;
		16'b0000001000010000 : data_out =  24'b000000000001010010110101;
		16'b0000001000010010 : data_out =  24'b000000000001010010111010;
		16'b0000001000010100 : data_out =  24'b000000000001010011000000;
		16'b0000001000010110 : data_out =  24'b000000000001010011000101;
		16'b0000001000011000 : data_out =  24'b000000000001010011001010;
		16'b0000001000011010 : data_out =  24'b000000000001010011010000;
		16'b0000001000011100 : data_out =  24'b000000000001010011010101;
		16'b0000001000011110 : data_out =  24'b000000000001010011011010;
		16'b0000001000100000 : data_out =  24'b000000000001010011100000;
		16'b0000001000100010 : data_out =  24'b000000000001010011100101;
		16'b0000001000100100 : data_out =  24'b000000000001010011101010;
		16'b0000001000100110 : data_out =  24'b000000000001010011110000;
		16'b0000001000101000 : data_out =  24'b000000000001010011110101;
		16'b0000001000101011 : data_out =  24'b000000000001010011111010;
		16'b0000001000101101 : data_out =  24'b000000000001010100000000;
		16'b0000001000101111 : data_out =  24'b000000000001010100000101;
		16'b0000001000110001 : data_out =  24'b000000000001010100001011;
		16'b0000001000110011 : data_out =  24'b000000000001010100010000;
		16'b0000001000110101 : data_out =  24'b000000000001010100010101;
		16'b0000001000110111 : data_out =  24'b000000000001010100011011;
		16'b0000001000111001 : data_out =  24'b000000000001010100100000;
		16'b0000001000111011 : data_out =  24'b000000000001010100100110;
		16'b0000001000111101 : data_out =  24'b000000000001010100101011;
		16'b0000001000111111 : data_out =  24'b000000000001010100110000;
		16'b0000001001000001 : data_out =  24'b000000000001010100110110;
		16'b0000001001000011 : data_out =  24'b000000000001010100111011;
		16'b0000001001000101 : data_out =  24'b000000000001010101000001;
		16'b0000001001000111 : data_out =  24'b000000000001010101000110;
		16'b0000001001001001 : data_out =  24'b000000000001010101001100;
		16'b0000001001001011 : data_out =  24'b000000000001010101010001;
		16'b0000001001001101 : data_out =  24'b000000000001010101010111;
		16'b0000001001001111 : data_out =  24'b000000000001010101011100;
		16'b0000001001010001 : data_out =  24'b000000000001010101100010;
		16'b0000001001010011 : data_out =  24'b000000000001010101100111;
		16'b0000001001010110 : data_out =  24'b000000000001010101101100;
		16'b0000001001011000 : data_out =  24'b000000000001010101110010;
		16'b0000001001011010 : data_out =  24'b000000000001010101110111;
		16'b0000001001011100 : data_out =  24'b000000000001010101111101;
		16'b0000001001011110 : data_out =  24'b000000000001010110000010;
		16'b0000001001100000 : data_out =  24'b000000000001010110001000;
		16'b0000001001100010 : data_out =  24'b000000000001010110001101;
		16'b0000001001100100 : data_out =  24'b000000000001010110010011;
		16'b0000001001100110 : data_out =  24'b000000000001010110011001;
		16'b0000001001101000 : data_out =  24'b000000000001010110011110;
		16'b0000001001101010 : data_out =  24'b000000000001010110100100;
		16'b0000001001101100 : data_out =  24'b000000000001010110101001;
		16'b0000001001101110 : data_out =  24'b000000000001010110101111;
		16'b0000001001110000 : data_out =  24'b000000000001010110110100;
		16'b0000001001110010 : data_out =  24'b000000000001010110111010;
		16'b0000001001110100 : data_out =  24'b000000000001010110111111;
		16'b0000001001110110 : data_out =  24'b000000000001010111000101;
		16'b0000001001111000 : data_out =  24'b000000000001010111001011;
		16'b0000001001111010 : data_out =  24'b000000000001010111010000;
		16'b0000001001111100 : data_out =  24'b000000000001010111010110;
		16'b0000001001111110 : data_out =  24'b000000000001010111011011;
		16'b0000001010000001 : data_out =  24'b000000000001010111100001;
		16'b0000001010000011 : data_out =  24'b000000000001010111100110;
		16'b0000001010000101 : data_out =  24'b000000000001010111101100;
		16'b0000001010000111 : data_out =  24'b000000000001010111110010;
		16'b0000001010001001 : data_out =  24'b000000000001010111110111;
		16'b0000001010001011 : data_out =  24'b000000000001010111111101;
		16'b0000001010001101 : data_out =  24'b000000000001011000000011;
		16'b0000001010001111 : data_out =  24'b000000000001011000001000;
		16'b0000001010010001 : data_out =  24'b000000000001011000001110;
		16'b0000001010010011 : data_out =  24'b000000000001011000010100;
		16'b0000001010010101 : data_out =  24'b000000000001011000011001;
		16'b0000001010010111 : data_out =  24'b000000000001011000011111;
		16'b0000001010011001 : data_out =  24'b000000000001011000100100;
		16'b0000001010011011 : data_out =  24'b000000000001011000101010;
		16'b0000001010011101 : data_out =  24'b000000000001011000110000;
		16'b0000001010011111 : data_out =  24'b000000000001011000110110;
		16'b0000001010100001 : data_out =  24'b000000000001011000111011;
		16'b0000001010100011 : data_out =  24'b000000000001011001000001;
		16'b0000001010100101 : data_out =  24'b000000000001011001000111;
		16'b0000001010100111 : data_out =  24'b000000000001011001001100;
		16'b0000001010101001 : data_out =  24'b000000000001011001010010;
		16'b0000001010101100 : data_out =  24'b000000000001011001011000;
		16'b0000001010101110 : data_out =  24'b000000000001011001011101;
		16'b0000001010110000 : data_out =  24'b000000000001011001100011;
		16'b0000001010110010 : data_out =  24'b000000000001011001101001;
		16'b0000001010110100 : data_out =  24'b000000000001011001101111;
		16'b0000001010110110 : data_out =  24'b000000000001011001110100;
		16'b0000001010111000 : data_out =  24'b000000000001011001111010;
		16'b0000001010111010 : data_out =  24'b000000000001011010000000;
		16'b0000001010111100 : data_out =  24'b000000000001011010000110;
		16'b0000001010111110 : data_out =  24'b000000000001011010001011;
		16'b0000001011000000 : data_out =  24'b000000000001011010010001;
		16'b0000001011000010 : data_out =  24'b000000000001011010010111;
		16'b0000001011000100 : data_out =  24'b000000000001011010011101;
		16'b0000001011000110 : data_out =  24'b000000000001011010100011;
		16'b0000001011001000 : data_out =  24'b000000000001011010101000;
		16'b0000001011001010 : data_out =  24'b000000000001011010101110;
		16'b0000001011001100 : data_out =  24'b000000000001011010110100;
		16'b0000001011001110 : data_out =  24'b000000000001011010111010;
		16'b0000001011010000 : data_out =  24'b000000000001011011000000;
		16'b0000001011010010 : data_out =  24'b000000000001011011000101;
		16'b0000001011010100 : data_out =  24'b000000000001011011001011;
		16'b0000001011010111 : data_out =  24'b000000000001011011010001;
		16'b0000001011011001 : data_out =  24'b000000000001011011010111;
		16'b0000001011011011 : data_out =  24'b000000000001011011011101;
		16'b0000001011011101 : data_out =  24'b000000000001011011100011;
		16'b0000001011011111 : data_out =  24'b000000000001011011101001;
		16'b0000001011100001 : data_out =  24'b000000000001011011101110;
		16'b0000001011100011 : data_out =  24'b000000000001011011110100;
		16'b0000001011100101 : data_out =  24'b000000000001011011111010;
		16'b0000001011100111 : data_out =  24'b000000000001011100000000;
		16'b0000001011101001 : data_out =  24'b000000000001011100000110;
		16'b0000001011101011 : data_out =  24'b000000000001011100001100;
		16'b0000001011101101 : data_out =  24'b000000000001011100010010;
		16'b0000001011101111 : data_out =  24'b000000000001011100011000;
		16'b0000001011110001 : data_out =  24'b000000000001011100011110;
		16'b0000001011110011 : data_out =  24'b000000000001011100100011;
		16'b0000001011110101 : data_out =  24'b000000000001011100101001;
		16'b0000001011110111 : data_out =  24'b000000000001011100101111;
		16'b0000001011111001 : data_out =  24'b000000000001011100110101;
		16'b0000001011111011 : data_out =  24'b000000000001011100111011;
		16'b0000001011111101 : data_out =  24'b000000000001011101000001;
		16'b0000001100000000 : data_out =  24'b000000000001011101000111;
		16'b0000001100000010 : data_out =  24'b000000000001011101001101;
		16'b0000001100000100 : data_out =  24'b000000000001011101010011;
		16'b0000001100000110 : data_out =  24'b000000000001011101011001;
		16'b0000001100001000 : data_out =  24'b000000000001011101011111;
		16'b0000001100001010 : data_out =  24'b000000000001011101100101;
		16'b0000001100001100 : data_out =  24'b000000000001011101101011;
		16'b0000001100001110 : data_out =  24'b000000000001011101110001;
		16'b0000001100010000 : data_out =  24'b000000000001011101110111;
		16'b0000001100010010 : data_out =  24'b000000000001011101111101;
		16'b0000001100010100 : data_out =  24'b000000000001011110000011;
		16'b0000001100010110 : data_out =  24'b000000000001011110001001;
		16'b0000001100011000 : data_out =  24'b000000000001011110001111;
		16'b0000001100011010 : data_out =  24'b000000000001011110010101;
		16'b0000001100011100 : data_out =  24'b000000000001011110011011;
		16'b0000001100011110 : data_out =  24'b000000000001011110100001;
		16'b0000001100100000 : data_out =  24'b000000000001011110100111;
		16'b0000001100100010 : data_out =  24'b000000000001011110101101;
		16'b0000001100100100 : data_out =  24'b000000000001011110110011;
		16'b0000001100100110 : data_out =  24'b000000000001011110111001;
		16'b0000001100101000 : data_out =  24'b000000000001011111000000;
		16'b0000001100101011 : data_out =  24'b000000000001011111000110;
		16'b0000001100101101 : data_out =  24'b000000000001011111001100;
		16'b0000001100101111 : data_out =  24'b000000000001011111010010;
		16'b0000001100110001 : data_out =  24'b000000000001011111011000;
		16'b0000001100110011 : data_out =  24'b000000000001011111011110;
		16'b0000001100110101 : data_out =  24'b000000000001011111100100;
		16'b0000001100110111 : data_out =  24'b000000000001011111101010;
		16'b0000001100111001 : data_out =  24'b000000000001011111110000;
		16'b0000001100111011 : data_out =  24'b000000000001011111110111;
		16'b0000001100111101 : data_out =  24'b000000000001011111111101;
		16'b0000001100111111 : data_out =  24'b000000000001100000000011;
		16'b0000001101000001 : data_out =  24'b000000000001100000001001;
		16'b0000001101000011 : data_out =  24'b000000000001100000001111;
		16'b0000001101000101 : data_out =  24'b000000000001100000010101;
		16'b0000001101000111 : data_out =  24'b000000000001100000011011;
		16'b0000001101001001 : data_out =  24'b000000000001100000100010;
		16'b0000001101001011 : data_out =  24'b000000000001100000101000;
		16'b0000001101001101 : data_out =  24'b000000000001100000101110;
		16'b0000001101001111 : data_out =  24'b000000000001100000110100;
		16'b0000001101010001 : data_out =  24'b000000000001100000111010;
		16'b0000001101010011 : data_out =  24'b000000000001100001000001;
		16'b0000001101010110 : data_out =  24'b000000000001100001000111;
		16'b0000001101011000 : data_out =  24'b000000000001100001001101;
		16'b0000001101011010 : data_out =  24'b000000000001100001010011;
		16'b0000001101011100 : data_out =  24'b000000000001100001011001;
		16'b0000001101011110 : data_out =  24'b000000000001100001100000;
		16'b0000001101100000 : data_out =  24'b000000000001100001100110;
		16'b0000001101100010 : data_out =  24'b000000000001100001101100;
		16'b0000001101100100 : data_out =  24'b000000000001100001110010;
		16'b0000001101100110 : data_out =  24'b000000000001100001111001;
		16'b0000001101101000 : data_out =  24'b000000000001100001111111;
		16'b0000001101101010 : data_out =  24'b000000000001100010000101;
		16'b0000001101101100 : data_out =  24'b000000000001100010001100;
		16'b0000001101101110 : data_out =  24'b000000000001100010010010;
		16'b0000001101110000 : data_out =  24'b000000000001100010011000;
		16'b0000001101110010 : data_out =  24'b000000000001100010011110;
		16'b0000001101110100 : data_out =  24'b000000000001100010100101;
		16'b0000001101110110 : data_out =  24'b000000000001100010101011;
		16'b0000001101111000 : data_out =  24'b000000000001100010110001;
		16'b0000001101111010 : data_out =  24'b000000000001100010111000;
		16'b0000001101111100 : data_out =  24'b000000000001100010111110;
		16'b0000001101111110 : data_out =  24'b000000000001100011000100;
		16'b0000001110000001 : data_out =  24'b000000000001100011001011;
		16'b0000001110000011 : data_out =  24'b000000000001100011010001;
		16'b0000001110000101 : data_out =  24'b000000000001100011010111;
		16'b0000001110000111 : data_out =  24'b000000000001100011011110;
		16'b0000001110001001 : data_out =  24'b000000000001100011100100;
		16'b0000001110001011 : data_out =  24'b000000000001100011101010;
		16'b0000001110001101 : data_out =  24'b000000000001100011110001;
		16'b0000001110001111 : data_out =  24'b000000000001100011110111;
		16'b0000001110010001 : data_out =  24'b000000000001100011111110;
		16'b0000001110010011 : data_out =  24'b000000000001100100000100;
		16'b0000001110010101 : data_out =  24'b000000000001100100001010;
		16'b0000001110010111 : data_out =  24'b000000000001100100010001;
		16'b0000001110011001 : data_out =  24'b000000000001100100010111;
		16'b0000001110011011 : data_out =  24'b000000000001100100011110;
		16'b0000001110011101 : data_out =  24'b000000000001100100100100;
		16'b0000001110011111 : data_out =  24'b000000000001100100101011;
		16'b0000001110100001 : data_out =  24'b000000000001100100110001;
		16'b0000001110100011 : data_out =  24'b000000000001100100111000;
		16'b0000001110100101 : data_out =  24'b000000000001100100111110;
		16'b0000001110100111 : data_out =  24'b000000000001100101000100;
		16'b0000001110101001 : data_out =  24'b000000000001100101001011;
		16'b0000001110101100 : data_out =  24'b000000000001100101010001;
		16'b0000001110101110 : data_out =  24'b000000000001100101011000;
		16'b0000001110110000 : data_out =  24'b000000000001100101011110;
		16'b0000001110110010 : data_out =  24'b000000000001100101100101;
		16'b0000001110110100 : data_out =  24'b000000000001100101101011;
		16'b0000001110110110 : data_out =  24'b000000000001100101110010;
		16'b0000001110111000 : data_out =  24'b000000000001100101111000;
		16'b0000001110111010 : data_out =  24'b000000000001100101111111;
		16'b0000001110111100 : data_out =  24'b000000000001100110000101;
		16'b0000001110111110 : data_out =  24'b000000000001100110001100;
		16'b0000001111000000 : data_out =  24'b000000000001100110010011;
		16'b0000001111000010 : data_out =  24'b000000000001100110011001;
		16'b0000001111000100 : data_out =  24'b000000000001100110100000;
		16'b0000001111000110 : data_out =  24'b000000000001100110100110;
		16'b0000001111001000 : data_out =  24'b000000000001100110101101;
		16'b0000001111001010 : data_out =  24'b000000000001100110110011;
		16'b0000001111001100 : data_out =  24'b000000000001100110111010;
		16'b0000001111001110 : data_out =  24'b000000000001100111000001;
		16'b0000001111010000 : data_out =  24'b000000000001100111000111;
		16'b0000001111010010 : data_out =  24'b000000000001100111001110;
		16'b0000001111010100 : data_out =  24'b000000000001100111010100;
		16'b0000001111010111 : data_out =  24'b000000000001100111011011;
		16'b0000001111011001 : data_out =  24'b000000000001100111100010;
		16'b0000001111011011 : data_out =  24'b000000000001100111101000;
		16'b0000001111011101 : data_out =  24'b000000000001100111101111;
		16'b0000001111011111 : data_out =  24'b000000000001100111110101;
		16'b0000001111100001 : data_out =  24'b000000000001100111111100;
		16'b0000001111100011 : data_out =  24'b000000000001101000000011;
		16'b0000001111100101 : data_out =  24'b000000000001101000001001;
		16'b0000001111100111 : data_out =  24'b000000000001101000010000;
		16'b0000001111101001 : data_out =  24'b000000000001101000010111;
		16'b0000001111101011 : data_out =  24'b000000000001101000011101;
		16'b0000001111101101 : data_out =  24'b000000000001101000100100;
		16'b0000001111101111 : data_out =  24'b000000000001101000101011;
		16'b0000001111110001 : data_out =  24'b000000000001101000110010;
		16'b0000001111110011 : data_out =  24'b000000000001101000111000;
		16'b0000001111110101 : data_out =  24'b000000000001101000111111;
		16'b0000001111110111 : data_out =  24'b000000000001101001000110;
		16'b0000001111111001 : data_out =  24'b000000000001101001001100;
		16'b0000001111111011 : data_out =  24'b000000000001101001010011;
		16'b0000001111111101 : data_out =  24'b000000000001101001011010;
		16'b0000010000000000 : data_out =  24'b000000000001101001100001;
		16'b0000010000000010 : data_out =  24'b000000000001101001100111;
		16'b0000010000000100 : data_out =  24'b000000000001101001101110;
		16'b0000010000000110 : data_out =  24'b000000000001101001110101;
		16'b0000010000001000 : data_out =  24'b000000000001101001111100;
		16'b0000010000001010 : data_out =  24'b000000000001101010000011;
		16'b0000010000001100 : data_out =  24'b000000000001101010001001;
		16'b0000010000001110 : data_out =  24'b000000000001101010010000;
		16'b0000010000010000 : data_out =  24'b000000000001101010010111;
		16'b0000010000010010 : data_out =  24'b000000000001101010011110;
		16'b0000010000010100 : data_out =  24'b000000000001101010100101;
		16'b0000010000010110 : data_out =  24'b000000000001101010101011;
		16'b0000010000011000 : data_out =  24'b000000000001101010110010;
		16'b0000010000011010 : data_out =  24'b000000000001101010111001;
		16'b0000010000011100 : data_out =  24'b000000000001101011000000;
		16'b0000010000011110 : data_out =  24'b000000000001101011000111;
		16'b0000010000100000 : data_out =  24'b000000000001101011001110;
		16'b0000010000100010 : data_out =  24'b000000000001101011010100;
		16'b0000010000100100 : data_out =  24'b000000000001101011011011;
		16'b0000010000100110 : data_out =  24'b000000000001101011100010;
		16'b0000010000101000 : data_out =  24'b000000000001101011101001;
		16'b0000010000101011 : data_out =  24'b000000000001101011110000;
		16'b0000010000101101 : data_out =  24'b000000000001101011110111;
		16'b0000010000101111 : data_out =  24'b000000000001101011111110;
		16'b0000010000110001 : data_out =  24'b000000000001101100000101;
		16'b0000010000110011 : data_out =  24'b000000000001101100001100;
		16'b0000010000110101 : data_out =  24'b000000000001101100010011;
		16'b0000010000110111 : data_out =  24'b000000000001101100011001;
		16'b0000010000111001 : data_out =  24'b000000000001101100100000;
		16'b0000010000111011 : data_out =  24'b000000000001101100100111;
		16'b0000010000111101 : data_out =  24'b000000000001101100101110;
		16'b0000010000111111 : data_out =  24'b000000000001101100110101;
		16'b0000010001000001 : data_out =  24'b000000000001101100111100;
		16'b0000010001000011 : data_out =  24'b000000000001101101000011;
		16'b0000010001000101 : data_out =  24'b000000000001101101001010;
		16'b0000010001000111 : data_out =  24'b000000000001101101010001;
		16'b0000010001001001 : data_out =  24'b000000000001101101011000;
		16'b0000010001001011 : data_out =  24'b000000000001101101011111;
		16'b0000010001001101 : data_out =  24'b000000000001101101100110;
		16'b0000010001001111 : data_out =  24'b000000000001101101101101;
		16'b0000010001010001 : data_out =  24'b000000000001101101110100;
		16'b0000010001010011 : data_out =  24'b000000000001101101111011;
		16'b0000010001010110 : data_out =  24'b000000000001101110000010;
		16'b0000010001011000 : data_out =  24'b000000000001101110001001;
		16'b0000010001011010 : data_out =  24'b000000000001101110010000;
		16'b0000010001011100 : data_out =  24'b000000000001101110010111;
		16'b0000010001011110 : data_out =  24'b000000000001101110011111;
		16'b0000010001100000 : data_out =  24'b000000000001101110100110;
		16'b0000010001100010 : data_out =  24'b000000000001101110101101;
		16'b0000010001100100 : data_out =  24'b000000000001101110110100;
		16'b0000010001100110 : data_out =  24'b000000000001101110111011;
		16'b0000010001101000 : data_out =  24'b000000000001101111000010;
		16'b0000010001101010 : data_out =  24'b000000000001101111001001;
		16'b0000010001101100 : data_out =  24'b000000000001101111010000;
		16'b0000010001101110 : data_out =  24'b000000000001101111010111;
		16'b0000010001110000 : data_out =  24'b000000000001101111011110;
		16'b0000010001110010 : data_out =  24'b000000000001101111100110;
		16'b0000010001110100 : data_out =  24'b000000000001101111101101;
		16'b0000010001110110 : data_out =  24'b000000000001101111110100;
		16'b0000010001111000 : data_out =  24'b000000000001101111111011;
		16'b0000010001111010 : data_out =  24'b000000000001110000000010;
		16'b0000010001111100 : data_out =  24'b000000000001110000001001;
		16'b0000010001111110 : data_out =  24'b000000000001110000010001;
		16'b0000010010000001 : data_out =  24'b000000000001110000011000;
		16'b0000010010000011 : data_out =  24'b000000000001110000011111;
		16'b0000010010000101 : data_out =  24'b000000000001110000100110;
		16'b0000010010000111 : data_out =  24'b000000000001110000101101;
		16'b0000010010001001 : data_out =  24'b000000000001110000110101;
		16'b0000010010001011 : data_out =  24'b000000000001110000111100;
		16'b0000010010001101 : data_out =  24'b000000000001110001000011;
		16'b0000010010001111 : data_out =  24'b000000000001110001001010;
		16'b0000010010010001 : data_out =  24'b000000000001110001010010;
		16'b0000010010010011 : data_out =  24'b000000000001110001011001;
		16'b0000010010010101 : data_out =  24'b000000000001110001100000;
		16'b0000010010010111 : data_out =  24'b000000000001110001100111;
		16'b0000010010011001 : data_out =  24'b000000000001110001101111;
		16'b0000010010011011 : data_out =  24'b000000000001110001110110;
		16'b0000010010011101 : data_out =  24'b000000000001110001111101;
		16'b0000010010011111 : data_out =  24'b000000000001110010000100;
		16'b0000010010100001 : data_out =  24'b000000000001110010001100;
		16'b0000010010100011 : data_out =  24'b000000000001110010010011;
		16'b0000010010100101 : data_out =  24'b000000000001110010011010;
		16'b0000010010100111 : data_out =  24'b000000000001110010100010;
		16'b0000010010101001 : data_out =  24'b000000000001110010101001;
		16'b0000010010101100 : data_out =  24'b000000000001110010110000;
		16'b0000010010101110 : data_out =  24'b000000000001110010111000;
		16'b0000010010110000 : data_out =  24'b000000000001110010111111;
		16'b0000010010110010 : data_out =  24'b000000000001110011000111;
		16'b0000010010110100 : data_out =  24'b000000000001110011001110;
		16'b0000010010110110 : data_out =  24'b000000000001110011010101;
		16'b0000010010111000 : data_out =  24'b000000000001110011011101;
		16'b0000010010111010 : data_out =  24'b000000000001110011100100;
		16'b0000010010111100 : data_out =  24'b000000000001110011101011;
		16'b0000010010111110 : data_out =  24'b000000000001110011110011;
		16'b0000010011000000 : data_out =  24'b000000000001110011111010;
		16'b0000010011000010 : data_out =  24'b000000000001110100000010;
		16'b0000010011000100 : data_out =  24'b000000000001110100001001;
		16'b0000010011000110 : data_out =  24'b000000000001110100010001;
		16'b0000010011001000 : data_out =  24'b000000000001110100011000;
		16'b0000010011001010 : data_out =  24'b000000000001110100011111;
		16'b0000010011001100 : data_out =  24'b000000000001110100100111;
		16'b0000010011001110 : data_out =  24'b000000000001110100101110;
		16'b0000010011010000 : data_out =  24'b000000000001110100110110;
		16'b0000010011010010 : data_out =  24'b000000000001110100111101;
		16'b0000010011010100 : data_out =  24'b000000000001110101000101;
		16'b0000010011010111 : data_out =  24'b000000000001110101001100;
		16'b0000010011011001 : data_out =  24'b000000000001110101010100;
		16'b0000010011011011 : data_out =  24'b000000000001110101011011;
		16'b0000010011011101 : data_out =  24'b000000000001110101100011;
		16'b0000010011011111 : data_out =  24'b000000000001110101101010;
		16'b0000010011100001 : data_out =  24'b000000000001110101110010;
		16'b0000010011100011 : data_out =  24'b000000000001110101111001;
		16'b0000010011100101 : data_out =  24'b000000000001110110000001;
		16'b0000010011100111 : data_out =  24'b000000000001110110001001;
		16'b0000010011101001 : data_out =  24'b000000000001110110010000;
		16'b0000010011101011 : data_out =  24'b000000000001110110011000;
		16'b0000010011101101 : data_out =  24'b000000000001110110011111;
		16'b0000010011101111 : data_out =  24'b000000000001110110100111;
		16'b0000010011110001 : data_out =  24'b000000000001110110101110;
		16'b0000010011110011 : data_out =  24'b000000000001110110110110;
		16'b0000010011110101 : data_out =  24'b000000000001110110111110;
		16'b0000010011110111 : data_out =  24'b000000000001110111000101;
		16'b0000010011111001 : data_out =  24'b000000000001110111001101;
		16'b0000010011111011 : data_out =  24'b000000000001110111010101;
		16'b0000010011111101 : data_out =  24'b000000000001110111011100;
		16'b0000010100000000 : data_out =  24'b000000000001110111100100;
		16'b0000010100000010 : data_out =  24'b000000000001110111101011;
		16'b0000010100000100 : data_out =  24'b000000000001110111110011;
		16'b0000010100000110 : data_out =  24'b000000000001110111111011;
		16'b0000010100001000 : data_out =  24'b000000000001111000000011;
		16'b0000010100001010 : data_out =  24'b000000000001111000001010;
		16'b0000010100001100 : data_out =  24'b000000000001111000010010;
		16'b0000010100001110 : data_out =  24'b000000000001111000011010;
		16'b0000010100010000 : data_out =  24'b000000000001111000100001;
		16'b0000010100010010 : data_out =  24'b000000000001111000101001;
		16'b0000010100010100 : data_out =  24'b000000000001111000110001;
		16'b0000010100010110 : data_out =  24'b000000000001111000111000;
		16'b0000010100011000 : data_out =  24'b000000000001111001000000;
		16'b0000010100011010 : data_out =  24'b000000000001111001001000;
		16'b0000010100011100 : data_out =  24'b000000000001111001010000;
		16'b0000010100011110 : data_out =  24'b000000000001111001010111;
		16'b0000010100100000 : data_out =  24'b000000000001111001011111;
		16'b0000010100100010 : data_out =  24'b000000000001111001100111;
		16'b0000010100100100 : data_out =  24'b000000000001111001101111;
		16'b0000010100100110 : data_out =  24'b000000000001111001110111;
		16'b0000010100101000 : data_out =  24'b000000000001111001111110;
		16'b0000010100101011 : data_out =  24'b000000000001111010000110;
		16'b0000010100101101 : data_out =  24'b000000000001111010001110;
		16'b0000010100101111 : data_out =  24'b000000000001111010010110;
		16'b0000010100110001 : data_out =  24'b000000000001111010011110;
		16'b0000010100110011 : data_out =  24'b000000000001111010100110;
		16'b0000010100110101 : data_out =  24'b000000000001111010101101;
		16'b0000010100110111 : data_out =  24'b000000000001111010110101;
		16'b0000010100111001 : data_out =  24'b000000000001111010111101;
		16'b0000010100111011 : data_out =  24'b000000000001111011000101;
		16'b0000010100111101 : data_out =  24'b000000000001111011001101;
		16'b0000010100111111 : data_out =  24'b000000000001111011010101;
		16'b0000010101000001 : data_out =  24'b000000000001111011011101;
		16'b0000010101000011 : data_out =  24'b000000000001111011100101;
		16'b0000010101000101 : data_out =  24'b000000000001111011101100;
		16'b0000010101000111 : data_out =  24'b000000000001111011110100;
		16'b0000010101001001 : data_out =  24'b000000000001111011111100;
		16'b0000010101001011 : data_out =  24'b000000000001111100000100;
		16'b0000010101001101 : data_out =  24'b000000000001111100001100;
		16'b0000010101001111 : data_out =  24'b000000000001111100010100;
		16'b0000010101010001 : data_out =  24'b000000000001111100011100;
		16'b0000010101010011 : data_out =  24'b000000000001111100100100;
		16'b0000010101010110 : data_out =  24'b000000000001111100101100;
		16'b0000010101011000 : data_out =  24'b000000000001111100110100;
		16'b0000010101011010 : data_out =  24'b000000000001111100111100;
		16'b0000010101011100 : data_out =  24'b000000000001111101000100;
		16'b0000010101011110 : data_out =  24'b000000000001111101001100;
		16'b0000010101100000 : data_out =  24'b000000000001111101010100;
		16'b0000010101100010 : data_out =  24'b000000000001111101011100;
		16'b0000010101100100 : data_out =  24'b000000000001111101100100;
		16'b0000010101100110 : data_out =  24'b000000000001111101101100;
		16'b0000010101101000 : data_out =  24'b000000000001111101110100;
		16'b0000010101101010 : data_out =  24'b000000000001111101111100;
		16'b0000010101101100 : data_out =  24'b000000000001111110000100;
		16'b0000010101101110 : data_out =  24'b000000000001111110001100;
		16'b0000010101110000 : data_out =  24'b000000000001111110010101;
		16'b0000010101110010 : data_out =  24'b000000000001111110011101;
		16'b0000010101110100 : data_out =  24'b000000000001111110100101;
		16'b0000010101110110 : data_out =  24'b000000000001111110101101;
		16'b0000010101111000 : data_out =  24'b000000000001111110110101;
		16'b0000010101111010 : data_out =  24'b000000000001111110111101;
		16'b0000010101111100 : data_out =  24'b000000000001111111000101;
		16'b0000010101111110 : data_out =  24'b000000000001111111001101;
		16'b0000010110000001 : data_out =  24'b000000000001111111010101;
		16'b0000010110000011 : data_out =  24'b000000000001111111011110;
		16'b0000010110000101 : data_out =  24'b000000000001111111100110;
		16'b0000010110000111 : data_out =  24'b000000000001111111101110;
		16'b0000010110001001 : data_out =  24'b000000000001111111110110;
		16'b0000010110001011 : data_out =  24'b000000000001111111111110;
		16'b0000010110001101 : data_out =  24'b000000000010000000000110;
		16'b0000010110001111 : data_out =  24'b000000000010000000001111;
		16'b0000010110010001 : data_out =  24'b000000000010000000010111;
		16'b0000010110010011 : data_out =  24'b000000000010000000011111;
		16'b0000010110010101 : data_out =  24'b000000000010000000100111;
		16'b0000010110010111 : data_out =  24'b000000000010000000110000;
		16'b0000010110011001 : data_out =  24'b000000000010000000111000;
		16'b0000010110011011 : data_out =  24'b000000000010000001000000;
		16'b0000010110011101 : data_out =  24'b000000000010000001001000;
		16'b0000010110011111 : data_out =  24'b000000000010000001010001;
		16'b0000010110100001 : data_out =  24'b000000000010000001011001;
		16'b0000010110100011 : data_out =  24'b000000000010000001100001;
		16'b0000010110100101 : data_out =  24'b000000000010000001101001;
		16'b0000010110100111 : data_out =  24'b000000000010000001110010;
		16'b0000010110101001 : data_out =  24'b000000000010000001111010;
		16'b0000010110101100 : data_out =  24'b000000000010000010000010;
		16'b0000010110101110 : data_out =  24'b000000000010000010001011;
		16'b0000010110110000 : data_out =  24'b000000000010000010010011;
		16'b0000010110110010 : data_out =  24'b000000000010000010011011;
		16'b0000010110110100 : data_out =  24'b000000000010000010100100;
		16'b0000010110110110 : data_out =  24'b000000000010000010101100;
		16'b0000010110111000 : data_out =  24'b000000000010000010110100;
		16'b0000010110111010 : data_out =  24'b000000000010000010111101;
		16'b0000010110111100 : data_out =  24'b000000000010000011000101;
		16'b0000010110111110 : data_out =  24'b000000000010000011001110;
		16'b0000010111000000 : data_out =  24'b000000000010000011010110;
		16'b0000010111000010 : data_out =  24'b000000000010000011011110;
		16'b0000010111000100 : data_out =  24'b000000000010000011100111;
		16'b0000010111000110 : data_out =  24'b000000000010000011101111;
		16'b0000010111001000 : data_out =  24'b000000000010000011111000;
		16'b0000010111001010 : data_out =  24'b000000000010000100000000;
		16'b0000010111001100 : data_out =  24'b000000000010000100001001;
		16'b0000010111001110 : data_out =  24'b000000000010000100010001;
		16'b0000010111010000 : data_out =  24'b000000000010000100011010;
		16'b0000010111010010 : data_out =  24'b000000000010000100100010;
		16'b0000010111010100 : data_out =  24'b000000000010000100101011;
		16'b0000010111010111 : data_out =  24'b000000000010000100110011;
		16'b0000010111011001 : data_out =  24'b000000000010000100111100;
		16'b0000010111011011 : data_out =  24'b000000000010000101000100;
		16'b0000010111011101 : data_out =  24'b000000000010000101001101;
		16'b0000010111011111 : data_out =  24'b000000000010000101010101;
		16'b0000010111100001 : data_out =  24'b000000000010000101011110;
		16'b0000010111100011 : data_out =  24'b000000000010000101100110;
		16'b0000010111100101 : data_out =  24'b000000000010000101101111;
		16'b0000010111100111 : data_out =  24'b000000000010000101110111;
		16'b0000010111101001 : data_out =  24'b000000000010000110000000;
		16'b0000010111101011 : data_out =  24'b000000000010000110001000;
		16'b0000010111101101 : data_out =  24'b000000000010000110010001;
		16'b0000010111101111 : data_out =  24'b000000000010000110011010;
		16'b0000010111110001 : data_out =  24'b000000000010000110100010;
		16'b0000010111110011 : data_out =  24'b000000000010000110101011;
		16'b0000010111110101 : data_out =  24'b000000000010000110110011;
		16'b0000010111110111 : data_out =  24'b000000000010000110111100;
		16'b0000010111111001 : data_out =  24'b000000000010000111000101;
		16'b0000010111111011 : data_out =  24'b000000000010000111001101;
		16'b0000010111111101 : data_out =  24'b000000000010000111010110;
		16'b0000011000000000 : data_out =  24'b000000000010000111011111;
		16'b0000011000000010 : data_out =  24'b000000000010000111100111;
		16'b0000011000000100 : data_out =  24'b000000000010000111110000;
		16'b0000011000000110 : data_out =  24'b000000000010000111111001;
		16'b0000011000001000 : data_out =  24'b000000000010001000000001;
		16'b0000011000001010 : data_out =  24'b000000000010001000001010;
		16'b0000011000001100 : data_out =  24'b000000000010001000010011;
		16'b0000011000001110 : data_out =  24'b000000000010001000011100;
		16'b0000011000010000 : data_out =  24'b000000000010001000100100;
		16'b0000011000010010 : data_out =  24'b000000000010001000101101;
		16'b0000011000010100 : data_out =  24'b000000000010001000110110;
		16'b0000011000010110 : data_out =  24'b000000000010001000111111;
		16'b0000011000011000 : data_out =  24'b000000000010001001000111;
		16'b0000011000011010 : data_out =  24'b000000000010001001010000;
		16'b0000011000011100 : data_out =  24'b000000000010001001011001;
		16'b0000011000011110 : data_out =  24'b000000000010001001100010;
		16'b0000011000100000 : data_out =  24'b000000000010001001101011;
		16'b0000011000100010 : data_out =  24'b000000000010001001110011;
		16'b0000011000100100 : data_out =  24'b000000000010001001111100;
		16'b0000011000100110 : data_out =  24'b000000000010001010000101;
		16'b0000011000101000 : data_out =  24'b000000000010001010001110;
		16'b0000011000101011 : data_out =  24'b000000000010001010010111;
		16'b0000011000101101 : data_out =  24'b000000000010001010100000;
		16'b0000011000101111 : data_out =  24'b000000000010001010101000;
		16'b0000011000110001 : data_out =  24'b000000000010001010110001;
		16'b0000011000110011 : data_out =  24'b000000000010001010111010;
		16'b0000011000110101 : data_out =  24'b000000000010001011000011;
		16'b0000011000110111 : data_out =  24'b000000000010001011001100;
		16'b0000011000111001 : data_out =  24'b000000000010001011010101;
		16'b0000011000111011 : data_out =  24'b000000000010001011011110;
		16'b0000011000111101 : data_out =  24'b000000000010001011100111;
		16'b0000011000111111 : data_out =  24'b000000000010001011110000;
		16'b0000011001000001 : data_out =  24'b000000000010001011111001;
		16'b0000011001000011 : data_out =  24'b000000000010001100000010;
		16'b0000011001000101 : data_out =  24'b000000000010001100001011;
		16'b0000011001000111 : data_out =  24'b000000000010001100010100;
		16'b0000011001001001 : data_out =  24'b000000000010001100011101;
		16'b0000011001001011 : data_out =  24'b000000000010001100100110;
		16'b0000011001001101 : data_out =  24'b000000000010001100101111;
		16'b0000011001001111 : data_out =  24'b000000000010001100111000;
		16'b0000011001010001 : data_out =  24'b000000000010001101000001;
		16'b0000011001010011 : data_out =  24'b000000000010001101001010;
		16'b0000011001010110 : data_out =  24'b000000000010001101010011;
		16'b0000011001011000 : data_out =  24'b000000000010001101011100;
		16'b0000011001011010 : data_out =  24'b000000000010001101100101;
		16'b0000011001011100 : data_out =  24'b000000000010001101101110;
		16'b0000011001011110 : data_out =  24'b000000000010001101110111;
		16'b0000011001100000 : data_out =  24'b000000000010001110000000;
		16'b0000011001100010 : data_out =  24'b000000000010001110001001;
		16'b0000011001100100 : data_out =  24'b000000000010001110010010;
		16'b0000011001100110 : data_out =  24'b000000000010001110011011;
		16'b0000011001101000 : data_out =  24'b000000000010001110100100;
		16'b0000011001101010 : data_out =  24'b000000000010001110101110;
		16'b0000011001101100 : data_out =  24'b000000000010001110110111;
		16'b0000011001101110 : data_out =  24'b000000000010001111000000;
		16'b0000011001110000 : data_out =  24'b000000000010001111001001;
		16'b0000011001110010 : data_out =  24'b000000000010001111010010;
		16'b0000011001110100 : data_out =  24'b000000000010001111011011;
		16'b0000011001110110 : data_out =  24'b000000000010001111100101;
		16'b0000011001111000 : data_out =  24'b000000000010001111101110;
		16'b0000011001111010 : data_out =  24'b000000000010001111110111;
		16'b0000011001111100 : data_out =  24'b000000000010010000000000;
		16'b0000011001111110 : data_out =  24'b000000000010010000001001;
		16'b0000011010000001 : data_out =  24'b000000000010010000010011;
		16'b0000011010000011 : data_out =  24'b000000000010010000011100;
		16'b0000011010000101 : data_out =  24'b000000000010010000100101;
		16'b0000011010000111 : data_out =  24'b000000000010010000101110;
		16'b0000011010001001 : data_out =  24'b000000000010010000111000;
		16'b0000011010001011 : data_out =  24'b000000000010010001000001;
		16'b0000011010001101 : data_out =  24'b000000000010010001001010;
		16'b0000011010001111 : data_out =  24'b000000000010010001010011;
		16'b0000011010010001 : data_out =  24'b000000000010010001011101;
		16'b0000011010010011 : data_out =  24'b000000000010010001100110;
		16'b0000011010010101 : data_out =  24'b000000000010010001101111;
		16'b0000011010010111 : data_out =  24'b000000000010010001111001;
		16'b0000011010011001 : data_out =  24'b000000000010010010000010;
		16'b0000011010011011 : data_out =  24'b000000000010010010001011;
		16'b0000011010011101 : data_out =  24'b000000000010010010010101;
		16'b0000011010011111 : data_out =  24'b000000000010010010011110;
		16'b0000011010100001 : data_out =  24'b000000000010010010101000;
		16'b0000011010100011 : data_out =  24'b000000000010010010110001;
		16'b0000011010100101 : data_out =  24'b000000000010010010111010;
		16'b0000011010100111 : data_out =  24'b000000000010010011000100;
		16'b0000011010101001 : data_out =  24'b000000000010010011001101;
		16'b0000011010101100 : data_out =  24'b000000000010010011010111;
		16'b0000011010101110 : data_out =  24'b000000000010010011100000;
		16'b0000011010110000 : data_out =  24'b000000000010010011101001;
		16'b0000011010110010 : data_out =  24'b000000000010010011110011;
		16'b0000011010110100 : data_out =  24'b000000000010010011111100;
		16'b0000011010110110 : data_out =  24'b000000000010010100000110;
		16'b0000011010111000 : data_out =  24'b000000000010010100001111;
		16'b0000011010111010 : data_out =  24'b000000000010010100011001;
		16'b0000011010111100 : data_out =  24'b000000000010010100100010;
		16'b0000011010111110 : data_out =  24'b000000000010010100101100;
		16'b0000011011000000 : data_out =  24'b000000000010010100110101;
		16'b0000011011000010 : data_out =  24'b000000000010010100111111;
		16'b0000011011000100 : data_out =  24'b000000000010010101001000;
		16'b0000011011000110 : data_out =  24'b000000000010010101010010;
		16'b0000011011001000 : data_out =  24'b000000000010010101011100;
		16'b0000011011001010 : data_out =  24'b000000000010010101100101;
		16'b0000011011001100 : data_out =  24'b000000000010010101101111;
		16'b0000011011001110 : data_out =  24'b000000000010010101111000;
		16'b0000011011010000 : data_out =  24'b000000000010010110000010;
		16'b0000011011010010 : data_out =  24'b000000000010010110001011;
		16'b0000011011010100 : data_out =  24'b000000000010010110010101;
		16'b0000011011010111 : data_out =  24'b000000000010010110011111;
		16'b0000011011011001 : data_out =  24'b000000000010010110101000;
		16'b0000011011011011 : data_out =  24'b000000000010010110110010;
		16'b0000011011011101 : data_out =  24'b000000000010010110111100;
		16'b0000011011011111 : data_out =  24'b000000000010010111000101;
		16'b0000011011100001 : data_out =  24'b000000000010010111001111;
		16'b0000011011100011 : data_out =  24'b000000000010010111011001;
		16'b0000011011100101 : data_out =  24'b000000000010010111100010;
		16'b0000011011100111 : data_out =  24'b000000000010010111101100;
		16'b0000011011101001 : data_out =  24'b000000000010010111110110;
		16'b0000011011101011 : data_out =  24'b000000000010011000000000;
		16'b0000011011101101 : data_out =  24'b000000000010011000001001;
		16'b0000011011101111 : data_out =  24'b000000000010011000010011;
		16'b0000011011110001 : data_out =  24'b000000000010011000011101;
		16'b0000011011110011 : data_out =  24'b000000000010011000100111;
		16'b0000011011110101 : data_out =  24'b000000000010011000110000;
		16'b0000011011110111 : data_out =  24'b000000000010011000111010;
		16'b0000011011111001 : data_out =  24'b000000000010011001000100;
		16'b0000011011111011 : data_out =  24'b000000000010011001001110;
		16'b0000011011111101 : data_out =  24'b000000000010011001010111;
		16'b0000011100000000 : data_out =  24'b000000000010011001100001;
		16'b0000011100000010 : data_out =  24'b000000000010011001101011;
		16'b0000011100000100 : data_out =  24'b000000000010011001110101;
		16'b0000011100000110 : data_out =  24'b000000000010011001111111;
		16'b0000011100001000 : data_out =  24'b000000000010011010001001;
		16'b0000011100001010 : data_out =  24'b000000000010011010010011;
		16'b0000011100001100 : data_out =  24'b000000000010011010011100;
		16'b0000011100001110 : data_out =  24'b000000000010011010100110;
		16'b0000011100010000 : data_out =  24'b000000000010011010110000;
		16'b0000011100010010 : data_out =  24'b000000000010011010111010;
		16'b0000011100010100 : data_out =  24'b000000000010011011000100;
		16'b0000011100010110 : data_out =  24'b000000000010011011001110;
		16'b0000011100011000 : data_out =  24'b000000000010011011011000;
		16'b0000011100011010 : data_out =  24'b000000000010011011100010;
		16'b0000011100011100 : data_out =  24'b000000000010011011101100;
		16'b0000011100011110 : data_out =  24'b000000000010011011110110;
		16'b0000011100100000 : data_out =  24'b000000000010011100000000;
		16'b0000011100100010 : data_out =  24'b000000000010011100001010;
		16'b0000011100100100 : data_out =  24'b000000000010011100010100;
		16'b0000011100100110 : data_out =  24'b000000000010011100011110;
		16'b0000011100101000 : data_out =  24'b000000000010011100101000;
		16'b0000011100101011 : data_out =  24'b000000000010011100110010;
		16'b0000011100101101 : data_out =  24'b000000000010011100111100;
		16'b0000011100101111 : data_out =  24'b000000000010011101000110;
		16'b0000011100110001 : data_out =  24'b000000000010011101010000;
		16'b0000011100110011 : data_out =  24'b000000000010011101011010;
		16'b0000011100110101 : data_out =  24'b000000000010011101100100;
		16'b0000011100110111 : data_out =  24'b000000000010011101101110;
		16'b0000011100111001 : data_out =  24'b000000000010011101111000;
		16'b0000011100111011 : data_out =  24'b000000000010011110000010;
		16'b0000011100111101 : data_out =  24'b000000000010011110001101;
		16'b0000011100111111 : data_out =  24'b000000000010011110010111;
		16'b0000011101000001 : data_out =  24'b000000000010011110100001;
		16'b0000011101000011 : data_out =  24'b000000000010011110101011;
		16'b0000011101000101 : data_out =  24'b000000000010011110110101;
		16'b0000011101000111 : data_out =  24'b000000000010011110111111;
		16'b0000011101001001 : data_out =  24'b000000000010011111001001;
		16'b0000011101001011 : data_out =  24'b000000000010011111010100;
		16'b0000011101001101 : data_out =  24'b000000000010011111011110;
		16'b0000011101001111 : data_out =  24'b000000000010011111101000;
		16'b0000011101010001 : data_out =  24'b000000000010011111110010;
		16'b0000011101010011 : data_out =  24'b000000000010011111111101;
		16'b0000011101010110 : data_out =  24'b000000000010100000000111;
		16'b0000011101011000 : data_out =  24'b000000000010100000010001;
		16'b0000011101011010 : data_out =  24'b000000000010100000011011;
		16'b0000011101011100 : data_out =  24'b000000000010100000100110;
		16'b0000011101011110 : data_out =  24'b000000000010100000110000;
		16'b0000011101100000 : data_out =  24'b000000000010100000111010;
		16'b0000011101100010 : data_out =  24'b000000000010100001000100;
		16'b0000011101100100 : data_out =  24'b000000000010100001001111;
		16'b0000011101100110 : data_out =  24'b000000000010100001011001;
		16'b0000011101101000 : data_out =  24'b000000000010100001100011;
		16'b0000011101101010 : data_out =  24'b000000000010100001101110;
		16'b0000011101101100 : data_out =  24'b000000000010100001111000;
		16'b0000011101101110 : data_out =  24'b000000000010100010000010;
		16'b0000011101110000 : data_out =  24'b000000000010100010001101;
		16'b0000011101110010 : data_out =  24'b000000000010100010010111;
		16'b0000011101110100 : data_out =  24'b000000000010100010100010;
		16'b0000011101110110 : data_out =  24'b000000000010100010101100;
		16'b0000011101111000 : data_out =  24'b000000000010100010110110;
		16'b0000011101111010 : data_out =  24'b000000000010100011000001;
		16'b0000011101111100 : data_out =  24'b000000000010100011001011;
		16'b0000011101111110 : data_out =  24'b000000000010100011010110;
		16'b0000011110000001 : data_out =  24'b000000000010100011100000;
		16'b0000011110000011 : data_out =  24'b000000000010100011101011;
		16'b0000011110000101 : data_out =  24'b000000000010100011110101;
		16'b0000011110000111 : data_out =  24'b000000000010100100000000;
		16'b0000011110001001 : data_out =  24'b000000000010100100001010;
		16'b0000011110001011 : data_out =  24'b000000000010100100010101;
		16'b0000011110001101 : data_out =  24'b000000000010100100011111;
		16'b0000011110001111 : data_out =  24'b000000000010100100101010;
		16'b0000011110010001 : data_out =  24'b000000000010100100110100;
		16'b0000011110010011 : data_out =  24'b000000000010100100111111;
		16'b0000011110010101 : data_out =  24'b000000000010100101001001;
		16'b0000011110010111 : data_out =  24'b000000000010100101010100;
		16'b0000011110011001 : data_out =  24'b000000000010100101011111;
		16'b0000011110011011 : data_out =  24'b000000000010100101101001;
		16'b0000011110011101 : data_out =  24'b000000000010100101110100;
		16'b0000011110011111 : data_out =  24'b000000000010100101111110;
		16'b0000011110100001 : data_out =  24'b000000000010100110001001;
		16'b0000011110100011 : data_out =  24'b000000000010100110010100;
		16'b0000011110100101 : data_out =  24'b000000000010100110011110;
		16'b0000011110100111 : data_out =  24'b000000000010100110101001;
		16'b0000011110101001 : data_out =  24'b000000000010100110110100;
		16'b0000011110101100 : data_out =  24'b000000000010100110111110;
		16'b0000011110101110 : data_out =  24'b000000000010100111001001;
		16'b0000011110110000 : data_out =  24'b000000000010100111010100;
		16'b0000011110110010 : data_out =  24'b000000000010100111011110;
		16'b0000011110110100 : data_out =  24'b000000000010100111101001;
		16'b0000011110110110 : data_out =  24'b000000000010100111110100;
		16'b0000011110111000 : data_out =  24'b000000000010100111111111;
		16'b0000011110111010 : data_out =  24'b000000000010101000001001;
		16'b0000011110111100 : data_out =  24'b000000000010101000010100;
		16'b0000011110111110 : data_out =  24'b000000000010101000011111;
		16'b0000011111000000 : data_out =  24'b000000000010101000101010;
		16'b0000011111000010 : data_out =  24'b000000000010101000110101;
		16'b0000011111000100 : data_out =  24'b000000000010101000111111;
		16'b0000011111000110 : data_out =  24'b000000000010101001001010;
		16'b0000011111001000 : data_out =  24'b000000000010101001010101;
		16'b0000011111001010 : data_out =  24'b000000000010101001100000;
		16'b0000011111001100 : data_out =  24'b000000000010101001101011;
		16'b0000011111001110 : data_out =  24'b000000000010101001110110;
		16'b0000011111010000 : data_out =  24'b000000000010101010000000;
		16'b0000011111010010 : data_out =  24'b000000000010101010001011;
		16'b0000011111010100 : data_out =  24'b000000000010101010010110;
		16'b0000011111010111 : data_out =  24'b000000000010101010100001;
		16'b0000011111011001 : data_out =  24'b000000000010101010101100;
		16'b0000011111011011 : data_out =  24'b000000000010101010110111;
		16'b0000011111011101 : data_out =  24'b000000000010101011000010;
		16'b0000011111011111 : data_out =  24'b000000000010101011001101;
		16'b0000011111100001 : data_out =  24'b000000000010101011011000;
		16'b0000011111100011 : data_out =  24'b000000000010101011100011;
		16'b0000011111100101 : data_out =  24'b000000000010101011101110;
		16'b0000011111100111 : data_out =  24'b000000000010101011111001;
		16'b0000011111101001 : data_out =  24'b000000000010101100000100;
		16'b0000011111101011 : data_out =  24'b000000000010101100001111;
		16'b0000011111101101 : data_out =  24'b000000000010101100011010;
		16'b0000011111101111 : data_out =  24'b000000000010101100100101;
		16'b0000011111110001 : data_out =  24'b000000000010101100110000;
		16'b0000011111110011 : data_out =  24'b000000000010101100111011;
		16'b0000011111110101 : data_out =  24'b000000000010101101000110;
		16'b0000011111110111 : data_out =  24'b000000000010101101010001;
		16'b0000011111111001 : data_out =  24'b000000000010101101011100;
		16'b0000011111111011 : data_out =  24'b000000000010101101100111;
		16'b0000011111111101 : data_out =  24'b000000000010101101110010;
		16'b0000100000000000 : data_out =  24'b000000000010101101111110;
		16'b0000100000000010 : data_out =  24'b000000000010101110001001;
		16'b0000100000000100 : data_out =  24'b000000000010101110010100;
		16'b0000100000000110 : data_out =  24'b000000000010101110011111;
		16'b0000100000001000 : data_out =  24'b000000000010101110101010;
		16'b0000100000001010 : data_out =  24'b000000000010101110110101;
		16'b0000100000001100 : data_out =  24'b000000000010101111000001;
		16'b0000100000001110 : data_out =  24'b000000000010101111001100;
		16'b0000100000010000 : data_out =  24'b000000000010101111010111;
		16'b0000100000010010 : data_out =  24'b000000000010101111100010;
		16'b0000100000010100 : data_out =  24'b000000000010101111101101;
		16'b0000100000010110 : data_out =  24'b000000000010101111111001;
		16'b0000100000011000 : data_out =  24'b000000000010110000000100;
		16'b0000100000011010 : data_out =  24'b000000000010110000001111;
		16'b0000100000011100 : data_out =  24'b000000000010110000011011;
		16'b0000100000011110 : data_out =  24'b000000000010110000100110;
		16'b0000100000100000 : data_out =  24'b000000000010110000110001;
		16'b0000100000100010 : data_out =  24'b000000000010110000111100;
		16'b0000100000100100 : data_out =  24'b000000000010110001001000;
		16'b0000100000100110 : data_out =  24'b000000000010110001010011;
		16'b0000100000101000 : data_out =  24'b000000000010110001011111;
		16'b0000100000101011 : data_out =  24'b000000000010110001101010;
		16'b0000100000101101 : data_out =  24'b000000000010110001110101;
		16'b0000100000101111 : data_out =  24'b000000000010110010000001;
		16'b0000100000110001 : data_out =  24'b000000000010110010001100;
		16'b0000100000110011 : data_out =  24'b000000000010110010010111;
		16'b0000100000110101 : data_out =  24'b000000000010110010100011;
		16'b0000100000110111 : data_out =  24'b000000000010110010101110;
		16'b0000100000111001 : data_out =  24'b000000000010110010111010;
		16'b0000100000111011 : data_out =  24'b000000000010110011000101;
		16'b0000100000111101 : data_out =  24'b000000000010110011010001;
		16'b0000100000111111 : data_out =  24'b000000000010110011011100;
		16'b0000100001000001 : data_out =  24'b000000000010110011101000;
		16'b0000100001000011 : data_out =  24'b000000000010110011110011;
		16'b0000100001000101 : data_out =  24'b000000000010110011111111;
		16'b0000100001000111 : data_out =  24'b000000000010110100001010;
		16'b0000100001001001 : data_out =  24'b000000000010110100010110;
		16'b0000100001001011 : data_out =  24'b000000000010110100100001;
		16'b0000100001001101 : data_out =  24'b000000000010110100101101;
		16'b0000100001001111 : data_out =  24'b000000000010110100111000;
		16'b0000100001010001 : data_out =  24'b000000000010110101000100;
		16'b0000100001010011 : data_out =  24'b000000000010110101010000;
		16'b0000100001010110 : data_out =  24'b000000000010110101011011;
		16'b0000100001011000 : data_out =  24'b000000000010110101100111;
		16'b0000100001011010 : data_out =  24'b000000000010110101110010;
		16'b0000100001011100 : data_out =  24'b000000000010110101111110;
		16'b0000100001011110 : data_out =  24'b000000000010110110001010;
		16'b0000100001100000 : data_out =  24'b000000000010110110010101;
		16'b0000100001100010 : data_out =  24'b000000000010110110100001;
		16'b0000100001100100 : data_out =  24'b000000000010110110101101;
		16'b0000100001100110 : data_out =  24'b000000000010110110111000;
		16'b0000100001101000 : data_out =  24'b000000000010110111000100;
		16'b0000100001101010 : data_out =  24'b000000000010110111010000;
		16'b0000100001101100 : data_out =  24'b000000000010110111011100;
		16'b0000100001101110 : data_out =  24'b000000000010110111100111;
		16'b0000100001110000 : data_out =  24'b000000000010110111110011;
		16'b0000100001110010 : data_out =  24'b000000000010110111111111;
		16'b0000100001110100 : data_out =  24'b000000000010111000001011;
		16'b0000100001110110 : data_out =  24'b000000000010111000010110;
		16'b0000100001111000 : data_out =  24'b000000000010111000100010;
		16'b0000100001111010 : data_out =  24'b000000000010111000101110;
		16'b0000100001111100 : data_out =  24'b000000000010111000111010;
		16'b0000100001111110 : data_out =  24'b000000000010111001000110;
		16'b0000100010000001 : data_out =  24'b000000000010111001010010;
		16'b0000100010000011 : data_out =  24'b000000000010111001011101;
		16'b0000100010000101 : data_out =  24'b000000000010111001101001;
		16'b0000100010000111 : data_out =  24'b000000000010111001110101;
		16'b0000100010001001 : data_out =  24'b000000000010111010000001;
		16'b0000100010001011 : data_out =  24'b000000000010111010001101;
		16'b0000100010001101 : data_out =  24'b000000000010111010011001;
		16'b0000100010001111 : data_out =  24'b000000000010111010100101;
		16'b0000100010010001 : data_out =  24'b000000000010111010110001;
		16'b0000100010010011 : data_out =  24'b000000000010111010111101;
		16'b0000100010010101 : data_out =  24'b000000000010111011001001;
		16'b0000100010010111 : data_out =  24'b000000000010111011010101;
		16'b0000100010011001 : data_out =  24'b000000000010111011100001;
		16'b0000100010011011 : data_out =  24'b000000000010111011101101;
		16'b0000100010011101 : data_out =  24'b000000000010111011111001;
		16'b0000100010011111 : data_out =  24'b000000000010111100000101;
		16'b0000100010100001 : data_out =  24'b000000000010111100010001;
		16'b0000100010100011 : data_out =  24'b000000000010111100011101;
		16'b0000100010100101 : data_out =  24'b000000000010111100101001;
		16'b0000100010100111 : data_out =  24'b000000000010111100110101;
		16'b0000100010101001 : data_out =  24'b000000000010111101000001;
		16'b0000100010101100 : data_out =  24'b000000000010111101001101;
		16'b0000100010101110 : data_out =  24'b000000000010111101011001;
		16'b0000100010110000 : data_out =  24'b000000000010111101100101;
		16'b0000100010110010 : data_out =  24'b000000000010111101110010;
		16'b0000100010110100 : data_out =  24'b000000000010111101111110;
		16'b0000100010110110 : data_out =  24'b000000000010111110001010;
		16'b0000100010111000 : data_out =  24'b000000000010111110010110;
		16'b0000100010111010 : data_out =  24'b000000000010111110100010;
		16'b0000100010111100 : data_out =  24'b000000000010111110101111;
		16'b0000100010111110 : data_out =  24'b000000000010111110111011;
		16'b0000100011000000 : data_out =  24'b000000000010111111000111;
		16'b0000100011000010 : data_out =  24'b000000000010111111010011;
		16'b0000100011000100 : data_out =  24'b000000000010111111011111;
		16'b0000100011000110 : data_out =  24'b000000000010111111101100;
		16'b0000100011001000 : data_out =  24'b000000000010111111111000;
		16'b0000100011001010 : data_out =  24'b000000000011000000000100;
		16'b0000100011001100 : data_out =  24'b000000000011000000010001;
		16'b0000100011001110 : data_out =  24'b000000000011000000011101;
		16'b0000100011010000 : data_out =  24'b000000000011000000101001;
		16'b0000100011010010 : data_out =  24'b000000000011000000110110;
		16'b0000100011010100 : data_out =  24'b000000000011000001000010;
		16'b0000100011010111 : data_out =  24'b000000000011000001001110;
		16'b0000100011011001 : data_out =  24'b000000000011000001011011;
		16'b0000100011011011 : data_out =  24'b000000000011000001100111;
		16'b0000100011011101 : data_out =  24'b000000000011000001110011;
		16'b0000100011011111 : data_out =  24'b000000000011000010000000;
		16'b0000100011100001 : data_out =  24'b000000000011000010001100;
		16'b0000100011100011 : data_out =  24'b000000000011000010011001;
		16'b0000100011100101 : data_out =  24'b000000000011000010100101;
		16'b0000100011100111 : data_out =  24'b000000000011000010110010;
		16'b0000100011101001 : data_out =  24'b000000000011000010111110;
		16'b0000100011101011 : data_out =  24'b000000000011000011001011;
		16'b0000100011101101 : data_out =  24'b000000000011000011010111;
		16'b0000100011101111 : data_out =  24'b000000000011000011100100;
		16'b0000100011110001 : data_out =  24'b000000000011000011110000;
		16'b0000100011110011 : data_out =  24'b000000000011000011111101;
		16'b0000100011110101 : data_out =  24'b000000000011000100001001;
		16'b0000100011110111 : data_out =  24'b000000000011000100010110;
		16'b0000100011111001 : data_out =  24'b000000000011000100100010;
		16'b0000100011111011 : data_out =  24'b000000000011000100101111;
		16'b0000100011111101 : data_out =  24'b000000000011000100111011;
		16'b0000100011111111 : data_out =  24'b000000000011000101001000;
		16'b0000100100000010 : data_out =  24'b000000000011000101010101;
		16'b0000100100000100 : data_out =  24'b000000000011000101100001;
		16'b0000100100000110 : data_out =  24'b000000000011000101101110;
		16'b0000100100001000 : data_out =  24'b000000000011000101111011;
		16'b0000100100001010 : data_out =  24'b000000000011000110000111;
		16'b0000100100001100 : data_out =  24'b000000000011000110010100;
		16'b0000100100001110 : data_out =  24'b000000000011000110100001;
		16'b0000100100010000 : data_out =  24'b000000000011000110101101;
		16'b0000100100010010 : data_out =  24'b000000000011000110111010;
		16'b0000100100010100 : data_out =  24'b000000000011000111000111;
		16'b0000100100010110 : data_out =  24'b000000000011000111010100;
		16'b0000100100011000 : data_out =  24'b000000000011000111100000;
		16'b0000100100011010 : data_out =  24'b000000000011000111101101;
		16'b0000100100011100 : data_out =  24'b000000000011000111111010;
		16'b0000100100011110 : data_out =  24'b000000000011001000000111;
		16'b0000100100100000 : data_out =  24'b000000000011001000010100;
		16'b0000100100100010 : data_out =  24'b000000000011001000100000;
		16'b0000100100100100 : data_out =  24'b000000000011001000101101;
		16'b0000100100100110 : data_out =  24'b000000000011001000111010;
		16'b0000100100101000 : data_out =  24'b000000000011001001000111;
		16'b0000100100101011 : data_out =  24'b000000000011001001010100;
		16'b0000100100101101 : data_out =  24'b000000000011001001100001;
		16'b0000100100101111 : data_out =  24'b000000000011001001101110;
		16'b0000100100110001 : data_out =  24'b000000000011001001111011;
		16'b0000100100110011 : data_out =  24'b000000000011001010000111;
		16'b0000100100110101 : data_out =  24'b000000000011001010010100;
		16'b0000100100110111 : data_out =  24'b000000000011001010100001;
		16'b0000100100111001 : data_out =  24'b000000000011001010101110;
		16'b0000100100111011 : data_out =  24'b000000000011001010111011;
		16'b0000100100111101 : data_out =  24'b000000000011001011001000;
		16'b0000100100111111 : data_out =  24'b000000000011001011010101;
		16'b0000100101000001 : data_out =  24'b000000000011001011100010;
		16'b0000100101000011 : data_out =  24'b000000000011001011101111;
		16'b0000100101000101 : data_out =  24'b000000000011001011111100;
		16'b0000100101000111 : data_out =  24'b000000000011001100001001;
		16'b0000100101001001 : data_out =  24'b000000000011001100010111;
		16'b0000100101001011 : data_out =  24'b000000000011001100100100;
		16'b0000100101001101 : data_out =  24'b000000000011001100110001;
		16'b0000100101001111 : data_out =  24'b000000000011001100111110;
		16'b0000100101010001 : data_out =  24'b000000000011001101001011;
		16'b0000100101010011 : data_out =  24'b000000000011001101011000;
		16'b0000100101010110 : data_out =  24'b000000000011001101100101;
		16'b0000100101011000 : data_out =  24'b000000000011001101110010;
		16'b0000100101011010 : data_out =  24'b000000000011001110000000;
		16'b0000100101011100 : data_out =  24'b000000000011001110001101;
		16'b0000100101011110 : data_out =  24'b000000000011001110011010;
		16'b0000100101100000 : data_out =  24'b000000000011001110100111;
		16'b0000100101100010 : data_out =  24'b000000000011001110110100;
		16'b0000100101100100 : data_out =  24'b000000000011001111000010;
		16'b0000100101100110 : data_out =  24'b000000000011001111001111;
		16'b0000100101101000 : data_out =  24'b000000000011001111011100;
		16'b0000100101101010 : data_out =  24'b000000000011001111101001;
		16'b0000100101101100 : data_out =  24'b000000000011001111110111;
		16'b0000100101101110 : data_out =  24'b000000000011010000000100;
		16'b0000100101110000 : data_out =  24'b000000000011010000010001;
		16'b0000100101110010 : data_out =  24'b000000000011010000011111;
		16'b0000100101110100 : data_out =  24'b000000000011010000101100;
		16'b0000100101110110 : data_out =  24'b000000000011010000111001;
		16'b0000100101111000 : data_out =  24'b000000000011010001000111;
		16'b0000100101111010 : data_out =  24'b000000000011010001010100;
		16'b0000100101111100 : data_out =  24'b000000000011010001100010;
		16'b0000100101111110 : data_out =  24'b000000000011010001101111;
		16'b0000100110000001 : data_out =  24'b000000000011010001111100;
		16'b0000100110000011 : data_out =  24'b000000000011010010001010;
		16'b0000100110000101 : data_out =  24'b000000000011010010010111;
		16'b0000100110000111 : data_out =  24'b000000000011010010100101;
		16'b0000100110001001 : data_out =  24'b000000000011010010110010;
		16'b0000100110001011 : data_out =  24'b000000000011010011000000;
		16'b0000100110001101 : data_out =  24'b000000000011010011001101;
		16'b0000100110001111 : data_out =  24'b000000000011010011011011;
		16'b0000100110010001 : data_out =  24'b000000000011010011101000;
		16'b0000100110010011 : data_out =  24'b000000000011010011110110;
		16'b0000100110010101 : data_out =  24'b000000000011010100000100;
		16'b0000100110010111 : data_out =  24'b000000000011010100010001;
		16'b0000100110011001 : data_out =  24'b000000000011010100011111;
		16'b0000100110011011 : data_out =  24'b000000000011010100101100;
		16'b0000100110011101 : data_out =  24'b000000000011010100111010;
		16'b0000100110011111 : data_out =  24'b000000000011010101001000;
		16'b0000100110100001 : data_out =  24'b000000000011010101010101;
		16'b0000100110100011 : data_out =  24'b000000000011010101100011;
		16'b0000100110100101 : data_out =  24'b000000000011010101110001;
		16'b0000100110100111 : data_out =  24'b000000000011010101111110;
		16'b0000100110101001 : data_out =  24'b000000000011010110001100;
		16'b0000100110101100 : data_out =  24'b000000000011010110011010;
		16'b0000100110101110 : data_out =  24'b000000000011010110100111;
		16'b0000100110110000 : data_out =  24'b000000000011010110110101;
		16'b0000100110110010 : data_out =  24'b000000000011010111000011;
		16'b0000100110110100 : data_out =  24'b000000000011010111010001;
		16'b0000100110110110 : data_out =  24'b000000000011010111011110;
		16'b0000100110111000 : data_out =  24'b000000000011010111101100;
		16'b0000100110111010 : data_out =  24'b000000000011010111111010;
		16'b0000100110111100 : data_out =  24'b000000000011011000001000;
		16'b0000100110111110 : data_out =  24'b000000000011011000010110;
		16'b0000100111000000 : data_out =  24'b000000000011011000100100;
		16'b0000100111000010 : data_out =  24'b000000000011011000110001;
		16'b0000100111000100 : data_out =  24'b000000000011011000111111;
		16'b0000100111000110 : data_out =  24'b000000000011011001001101;
		16'b0000100111001000 : data_out =  24'b000000000011011001011011;
		16'b0000100111001010 : data_out =  24'b000000000011011001101001;
		16'b0000100111001100 : data_out =  24'b000000000011011001110111;
		16'b0000100111001110 : data_out =  24'b000000000011011010000101;
		16'b0000100111010000 : data_out =  24'b000000000011011010010011;
		16'b0000100111010010 : data_out =  24'b000000000011011010100001;
		16'b0000100111010100 : data_out =  24'b000000000011011010101111;
		16'b0000100111010111 : data_out =  24'b000000000011011010111101;
		16'b0000100111011001 : data_out =  24'b000000000011011011001011;
		16'b0000100111011011 : data_out =  24'b000000000011011011011001;
		16'b0000100111011101 : data_out =  24'b000000000011011011100111;
		16'b0000100111011111 : data_out =  24'b000000000011011011110101;
		16'b0000100111100001 : data_out =  24'b000000000011011100000011;
		16'b0000100111100011 : data_out =  24'b000000000011011100010001;
		16'b0000100111100101 : data_out =  24'b000000000011011100011111;
		16'b0000100111100111 : data_out =  24'b000000000011011100101101;
		16'b0000100111101001 : data_out =  24'b000000000011011100111100;
		16'b0000100111101011 : data_out =  24'b000000000011011101001010;
		16'b0000100111101101 : data_out =  24'b000000000011011101011000;
		16'b0000100111101111 : data_out =  24'b000000000011011101100110;
		16'b0000100111110001 : data_out =  24'b000000000011011101110100;
		16'b0000100111110011 : data_out =  24'b000000000011011110000010;
		16'b0000100111110101 : data_out =  24'b000000000011011110010001;
		16'b0000100111110111 : data_out =  24'b000000000011011110011111;
		16'b0000100111111001 : data_out =  24'b000000000011011110101101;
		16'b0000100111111011 : data_out =  24'b000000000011011110111011;
		16'b0000100111111101 : data_out =  24'b000000000011011111001010;
		16'b0000100111111111 : data_out =  24'b000000000011011111011000;
		16'b0000101000000010 : data_out =  24'b000000000011011111100110;
		16'b0000101000000100 : data_out =  24'b000000000011011111110101;
		16'b0000101000000110 : data_out =  24'b000000000011100000000011;
		16'b0000101000001000 : data_out =  24'b000000000011100000010001;
		16'b0000101000001010 : data_out =  24'b000000000011100000100000;
		16'b0000101000001100 : data_out =  24'b000000000011100000101110;
		16'b0000101000001110 : data_out =  24'b000000000011100000111100;
		16'b0000101000010000 : data_out =  24'b000000000011100001001011;
		16'b0000101000010010 : data_out =  24'b000000000011100001011001;
		16'b0000101000010100 : data_out =  24'b000000000011100001101000;
		16'b0000101000010110 : data_out =  24'b000000000011100001110110;
		16'b0000101000011000 : data_out =  24'b000000000011100010000101;
		16'b0000101000011010 : data_out =  24'b000000000011100010010011;
		16'b0000101000011100 : data_out =  24'b000000000011100010100010;
		16'b0000101000011110 : data_out =  24'b000000000011100010110000;
		16'b0000101000100000 : data_out =  24'b000000000011100010111111;
		16'b0000101000100010 : data_out =  24'b000000000011100011001101;
		16'b0000101000100100 : data_out =  24'b000000000011100011011100;
		16'b0000101000100110 : data_out =  24'b000000000011100011101010;
		16'b0000101000101000 : data_out =  24'b000000000011100011111001;
		16'b0000101000101011 : data_out =  24'b000000000011100100000111;
		16'b0000101000101101 : data_out =  24'b000000000011100100010110;
		16'b0000101000101111 : data_out =  24'b000000000011100100100101;
		16'b0000101000110001 : data_out =  24'b000000000011100100110011;
		16'b0000101000110011 : data_out =  24'b000000000011100101000010;
		16'b0000101000110101 : data_out =  24'b000000000011100101010001;
		16'b0000101000110111 : data_out =  24'b000000000011100101011111;
		16'b0000101000111001 : data_out =  24'b000000000011100101101110;
		16'b0000101000111011 : data_out =  24'b000000000011100101111101;
		16'b0000101000111101 : data_out =  24'b000000000011100110001011;
		16'b0000101000111111 : data_out =  24'b000000000011100110011010;
		16'b0000101001000001 : data_out =  24'b000000000011100110101001;
		16'b0000101001000011 : data_out =  24'b000000000011100110111000;
		16'b0000101001000101 : data_out =  24'b000000000011100111000110;
		16'b0000101001000111 : data_out =  24'b000000000011100111010101;
		16'b0000101001001001 : data_out =  24'b000000000011100111100100;
		16'b0000101001001011 : data_out =  24'b000000000011100111110011;
		16'b0000101001001101 : data_out =  24'b000000000011101000000010;
		16'b0000101001001111 : data_out =  24'b000000000011101000010001;
		16'b0000101001010001 : data_out =  24'b000000000011101000011111;
		16'b0000101001010011 : data_out =  24'b000000000011101000101110;
		16'b0000101001010110 : data_out =  24'b000000000011101000111101;
		16'b0000101001011000 : data_out =  24'b000000000011101001001100;
		16'b0000101001011010 : data_out =  24'b000000000011101001011011;
		16'b0000101001011100 : data_out =  24'b000000000011101001101010;
		16'b0000101001011110 : data_out =  24'b000000000011101001111001;
		16'b0000101001100000 : data_out =  24'b000000000011101010001000;
		16'b0000101001100010 : data_out =  24'b000000000011101010010111;
		16'b0000101001100100 : data_out =  24'b000000000011101010100110;
		16'b0000101001100110 : data_out =  24'b000000000011101010110101;
		16'b0000101001101000 : data_out =  24'b000000000011101011000100;
		16'b0000101001101010 : data_out =  24'b000000000011101011010011;
		16'b0000101001101100 : data_out =  24'b000000000011101011100010;
		16'b0000101001101110 : data_out =  24'b000000000011101011110001;
		16'b0000101001110000 : data_out =  24'b000000000011101100000000;
		16'b0000101001110010 : data_out =  24'b000000000011101100001111;
		16'b0000101001110100 : data_out =  24'b000000000011101100011111;
		16'b0000101001110110 : data_out =  24'b000000000011101100101110;
		16'b0000101001111000 : data_out =  24'b000000000011101100111101;
		16'b0000101001111010 : data_out =  24'b000000000011101101001100;
		16'b0000101001111100 : data_out =  24'b000000000011101101011011;
		16'b0000101001111110 : data_out =  24'b000000000011101101101010;
		16'b0000101010000001 : data_out =  24'b000000000011101101111010;
		16'b0000101010000011 : data_out =  24'b000000000011101110001001;
		16'b0000101010000101 : data_out =  24'b000000000011101110011000;
		16'b0000101010000111 : data_out =  24'b000000000011101110100111;
		16'b0000101010001001 : data_out =  24'b000000000011101110110111;
		16'b0000101010001011 : data_out =  24'b000000000011101111000110;
		16'b0000101010001101 : data_out =  24'b000000000011101111010101;
		16'b0000101010001111 : data_out =  24'b000000000011101111100101;
		16'b0000101010010001 : data_out =  24'b000000000011101111110100;
		16'b0000101010010011 : data_out =  24'b000000000011110000000011;
		16'b0000101010010101 : data_out =  24'b000000000011110000010011;
		16'b0000101010010111 : data_out =  24'b000000000011110000100010;
		16'b0000101010011001 : data_out =  24'b000000000011110000110001;
		16'b0000101010011011 : data_out =  24'b000000000011110001000001;
		16'b0000101010011101 : data_out =  24'b000000000011110001010000;
		16'b0000101010011111 : data_out =  24'b000000000011110001100000;
		16'b0000101010100001 : data_out =  24'b000000000011110001101111;
		16'b0000101010100011 : data_out =  24'b000000000011110001111111;
		16'b0000101010100101 : data_out =  24'b000000000011110010001110;
		16'b0000101010100111 : data_out =  24'b000000000011110010011110;
		16'b0000101010101001 : data_out =  24'b000000000011110010101101;
		16'b0000101010101100 : data_out =  24'b000000000011110010111101;
		16'b0000101010101110 : data_out =  24'b000000000011110011001100;
		16'b0000101010110000 : data_out =  24'b000000000011110011011100;
		16'b0000101010110010 : data_out =  24'b000000000011110011101011;
		16'b0000101010110100 : data_out =  24'b000000000011110011111011;
		16'b0000101010110110 : data_out =  24'b000000000011110100001011;
		16'b0000101010111000 : data_out =  24'b000000000011110100011010;
		16'b0000101010111010 : data_out =  24'b000000000011110100101010;
		16'b0000101010111100 : data_out =  24'b000000000011110100111010;
		16'b0000101010111110 : data_out =  24'b000000000011110101001001;
		16'b0000101011000000 : data_out =  24'b000000000011110101011001;
		16'b0000101011000010 : data_out =  24'b000000000011110101101001;
		16'b0000101011000100 : data_out =  24'b000000000011110101111000;
		16'b0000101011000110 : data_out =  24'b000000000011110110001000;
		16'b0000101011001000 : data_out =  24'b000000000011110110011000;
		16'b0000101011001010 : data_out =  24'b000000000011110110101000;
		16'b0000101011001100 : data_out =  24'b000000000011110110111000;
		16'b0000101011001110 : data_out =  24'b000000000011110111000111;
		16'b0000101011010000 : data_out =  24'b000000000011110111010111;
		16'b0000101011010010 : data_out =  24'b000000000011110111100111;
		16'b0000101011010100 : data_out =  24'b000000000011110111110111;
		16'b0000101011010111 : data_out =  24'b000000000011111000000111;
		16'b0000101011011001 : data_out =  24'b000000000011111000010111;
		16'b0000101011011011 : data_out =  24'b000000000011111000100111;
		16'b0000101011011101 : data_out =  24'b000000000011111000110110;
		16'b0000101011011111 : data_out =  24'b000000000011111001000110;
		16'b0000101011100001 : data_out =  24'b000000000011111001010110;
		16'b0000101011100011 : data_out =  24'b000000000011111001100110;
		16'b0000101011100101 : data_out =  24'b000000000011111001110110;
		16'b0000101011100111 : data_out =  24'b000000000011111010000110;
		16'b0000101011101001 : data_out =  24'b000000000011111010010110;
		16'b0000101011101011 : data_out =  24'b000000000011111010100110;
		16'b0000101011101101 : data_out =  24'b000000000011111010110110;
		16'b0000101011101111 : data_out =  24'b000000000011111011000110;
		16'b0000101011110001 : data_out =  24'b000000000011111011010110;
		16'b0000101011110011 : data_out =  24'b000000000011111011100111;
		16'b0000101011110101 : data_out =  24'b000000000011111011110111;
		16'b0000101011110111 : data_out =  24'b000000000011111100000111;
		16'b0000101011111001 : data_out =  24'b000000000011111100010111;
		16'b0000101011111011 : data_out =  24'b000000000011111100100111;
		16'b0000101011111101 : data_out =  24'b000000000011111100110111;
		16'b0000101011111111 : data_out =  24'b000000000011111101000111;
		16'b0000101100000010 : data_out =  24'b000000000011111101011000;
		16'b0000101100000100 : data_out =  24'b000000000011111101101000;
		16'b0000101100000110 : data_out =  24'b000000000011111101111000;
		16'b0000101100001000 : data_out =  24'b000000000011111110001000;
		16'b0000101100001010 : data_out =  24'b000000000011111110011001;
		16'b0000101100001100 : data_out =  24'b000000000011111110101001;
		16'b0000101100001110 : data_out =  24'b000000000011111110111001;
		16'b0000101100010000 : data_out =  24'b000000000011111111001010;
		16'b0000101100010010 : data_out =  24'b000000000011111111011010;
		16'b0000101100010100 : data_out =  24'b000000000011111111101010;
		16'b0000101100010110 : data_out =  24'b000000000011111111111011;
		16'b0000101100011000 : data_out =  24'b000000000100000000001011;
		16'b0000101100011010 : data_out =  24'b000000000100000000011011;
		16'b0000101100011100 : data_out =  24'b000000000100000000101100;
		16'b0000101100011110 : data_out =  24'b000000000100000000111100;
		16'b0000101100100000 : data_out =  24'b000000000100000001001101;
		16'b0000101100100010 : data_out =  24'b000000000100000001011101;
		16'b0000101100100100 : data_out =  24'b000000000100000001101110;
		16'b0000101100100110 : data_out =  24'b000000000100000001111110;
		16'b0000101100101000 : data_out =  24'b000000000100000010001111;
		16'b0000101100101011 : data_out =  24'b000000000100000010011111;
		16'b0000101100101101 : data_out =  24'b000000000100000010110000;
		16'b0000101100101111 : data_out =  24'b000000000100000011000000;
		16'b0000101100110001 : data_out =  24'b000000000100000011010001;
		16'b0000101100110011 : data_out =  24'b000000000100000011100010;
		16'b0000101100110101 : data_out =  24'b000000000100000011110010;
		16'b0000101100110111 : data_out =  24'b000000000100000100000011;
		16'b0000101100111001 : data_out =  24'b000000000100000100010100;
		16'b0000101100111011 : data_out =  24'b000000000100000100100100;
		16'b0000101100111101 : data_out =  24'b000000000100000100110101;
		16'b0000101100111111 : data_out =  24'b000000000100000101000110;
		16'b0000101101000001 : data_out =  24'b000000000100000101010110;
		16'b0000101101000011 : data_out =  24'b000000000100000101100111;
		16'b0000101101000101 : data_out =  24'b000000000100000101111000;
		16'b0000101101000111 : data_out =  24'b000000000100000110001001;
		16'b0000101101001001 : data_out =  24'b000000000100000110011001;
		16'b0000101101001011 : data_out =  24'b000000000100000110101010;
		16'b0000101101001101 : data_out =  24'b000000000100000110111011;
		16'b0000101101001111 : data_out =  24'b000000000100000111001100;
		16'b0000101101010001 : data_out =  24'b000000000100000111011101;
		16'b0000101101010011 : data_out =  24'b000000000100000111101101;
		16'b0000101101010110 : data_out =  24'b000000000100000111111110;
		16'b0000101101011000 : data_out =  24'b000000000100001000001111;
		16'b0000101101011010 : data_out =  24'b000000000100001000100000;
		16'b0000101101011100 : data_out =  24'b000000000100001000110001;
		16'b0000101101011110 : data_out =  24'b000000000100001001000010;
		16'b0000101101100000 : data_out =  24'b000000000100001001010011;
		16'b0000101101100010 : data_out =  24'b000000000100001001100100;
		16'b0000101101100100 : data_out =  24'b000000000100001001110101;
		16'b0000101101100110 : data_out =  24'b000000000100001010000110;
		16'b0000101101101000 : data_out =  24'b000000000100001010010111;
		16'b0000101101101010 : data_out =  24'b000000000100001010101000;
		16'b0000101101101100 : data_out =  24'b000000000100001010111001;
		16'b0000101101101110 : data_out =  24'b000000000100001011001010;
		16'b0000101101110000 : data_out =  24'b000000000100001011011011;
		16'b0000101101110010 : data_out =  24'b000000000100001011101101;
		16'b0000101101110100 : data_out =  24'b000000000100001011111110;
		16'b0000101101110110 : data_out =  24'b000000000100001100001111;
		16'b0000101101111000 : data_out =  24'b000000000100001100100000;
		16'b0000101101111010 : data_out =  24'b000000000100001100110001;
		16'b0000101101111100 : data_out =  24'b000000000100001101000010;
		16'b0000101101111110 : data_out =  24'b000000000100001101010100;
		16'b0000101110000001 : data_out =  24'b000000000100001101100101;
		16'b0000101110000011 : data_out =  24'b000000000100001101110110;
		16'b0000101110000101 : data_out =  24'b000000000100001110000111;
		16'b0000101110000111 : data_out =  24'b000000000100001110011001;
		16'b0000101110001001 : data_out =  24'b000000000100001110101010;
		16'b0000101110001011 : data_out =  24'b000000000100001110111011;
		16'b0000101110001101 : data_out =  24'b000000000100001111001101;
		16'b0000101110001111 : data_out =  24'b000000000100001111011110;
		16'b0000101110010001 : data_out =  24'b000000000100001111110000;
		16'b0000101110010011 : data_out =  24'b000000000100010000000001;
		16'b0000101110010101 : data_out =  24'b000000000100010000010010;
		16'b0000101110010111 : data_out =  24'b000000000100010000100100;
		16'b0000101110011001 : data_out =  24'b000000000100010000110101;
		16'b0000101110011011 : data_out =  24'b000000000100010001000111;
		16'b0000101110011101 : data_out =  24'b000000000100010001011000;
		16'b0000101110011111 : data_out =  24'b000000000100010001101010;
		16'b0000101110100001 : data_out =  24'b000000000100010001111011;
		16'b0000101110100011 : data_out =  24'b000000000100010010001101;
		16'b0000101110100101 : data_out =  24'b000000000100010010011110;
		16'b0000101110100111 : data_out =  24'b000000000100010010110000;
		16'b0000101110101001 : data_out =  24'b000000000100010011000001;
		16'b0000101110101100 : data_out =  24'b000000000100010011010011;
		16'b0000101110101110 : data_out =  24'b000000000100010011100101;
		16'b0000101110110000 : data_out =  24'b000000000100010011110110;
		16'b0000101110110010 : data_out =  24'b000000000100010100001000;
		16'b0000101110110100 : data_out =  24'b000000000100010100011010;
		16'b0000101110110110 : data_out =  24'b000000000100010100101011;
		16'b0000101110111000 : data_out =  24'b000000000100010100111101;
		16'b0000101110111010 : data_out =  24'b000000000100010101001111;
		16'b0000101110111100 : data_out =  24'b000000000100010101100001;
		16'b0000101110111110 : data_out =  24'b000000000100010101110010;
		16'b0000101111000000 : data_out =  24'b000000000100010110000100;
		16'b0000101111000010 : data_out =  24'b000000000100010110010110;
		16'b0000101111000100 : data_out =  24'b000000000100010110101000;
		16'b0000101111000110 : data_out =  24'b000000000100010110111010;
		16'b0000101111001000 : data_out =  24'b000000000100010111001011;
		16'b0000101111001010 : data_out =  24'b000000000100010111011101;
		16'b0000101111001100 : data_out =  24'b000000000100010111101111;
		16'b0000101111001110 : data_out =  24'b000000000100011000000001;
		16'b0000101111010000 : data_out =  24'b000000000100011000010011;
		16'b0000101111010010 : data_out =  24'b000000000100011000100101;
		16'b0000101111010100 : data_out =  24'b000000000100011000110111;
		16'b0000101111010111 : data_out =  24'b000000000100011001001001;
		16'b0000101111011001 : data_out =  24'b000000000100011001011011;
		16'b0000101111011011 : data_out =  24'b000000000100011001101101;
		16'b0000101111011101 : data_out =  24'b000000000100011001111111;
		16'b0000101111011111 : data_out =  24'b000000000100011010010001;
		16'b0000101111100001 : data_out =  24'b000000000100011010100011;
		16'b0000101111100011 : data_out =  24'b000000000100011010110101;
		16'b0000101111100101 : data_out =  24'b000000000100011011000111;
		16'b0000101111100111 : data_out =  24'b000000000100011011011010;
		16'b0000101111101001 : data_out =  24'b000000000100011011101100;
		16'b0000101111101011 : data_out =  24'b000000000100011011111110;
		16'b0000101111101101 : data_out =  24'b000000000100011100010000;
		16'b0000101111101111 : data_out =  24'b000000000100011100100010;
		16'b0000101111110001 : data_out =  24'b000000000100011100110100;
		16'b0000101111110011 : data_out =  24'b000000000100011101000111;
		16'b0000101111110101 : data_out =  24'b000000000100011101011001;
		16'b0000101111110111 : data_out =  24'b000000000100011101101011;
		16'b0000101111111001 : data_out =  24'b000000000100011101111110;
		16'b0000101111111011 : data_out =  24'b000000000100011110010000;
		16'b0000101111111101 : data_out =  24'b000000000100011110100010;
		16'b0000101111111111 : data_out =  24'b000000000100011110110100;
		16'b0000110000000010 : data_out =  24'b000000000100011111000111;
		16'b0000110000000100 : data_out =  24'b000000000100011111011001;
		16'b0000110000000110 : data_out =  24'b000000000100011111101100;
		16'b0000110000001000 : data_out =  24'b000000000100011111111110;
		16'b0000110000001010 : data_out =  24'b000000000100100000010001;
		16'b0000110000001100 : data_out =  24'b000000000100100000100011;
		16'b0000110000001110 : data_out =  24'b000000000100100000110101;
		16'b0000110000010000 : data_out =  24'b000000000100100001001000;
		16'b0000110000010010 : data_out =  24'b000000000100100001011010;
		16'b0000110000010100 : data_out =  24'b000000000100100001101101;
		16'b0000110000010110 : data_out =  24'b000000000100100010000000;
		16'b0000110000011000 : data_out =  24'b000000000100100010010010;
		16'b0000110000011010 : data_out =  24'b000000000100100010100101;
		16'b0000110000011100 : data_out =  24'b000000000100100010110111;
		16'b0000110000011110 : data_out =  24'b000000000100100011001010;
		16'b0000110000100000 : data_out =  24'b000000000100100011011101;
		16'b0000110000100010 : data_out =  24'b000000000100100011101111;
		16'b0000110000100100 : data_out =  24'b000000000100100100000010;
		16'b0000110000100110 : data_out =  24'b000000000100100100010101;
		16'b0000110000101000 : data_out =  24'b000000000100100100100111;
		16'b0000110000101011 : data_out =  24'b000000000100100100111010;
		16'b0000110000101101 : data_out =  24'b000000000100100101001101;
		16'b0000110000101111 : data_out =  24'b000000000100100101100000;
		16'b0000110000110001 : data_out =  24'b000000000100100101110010;
		16'b0000110000110011 : data_out =  24'b000000000100100110000101;
		16'b0000110000110101 : data_out =  24'b000000000100100110011000;
		16'b0000110000110111 : data_out =  24'b000000000100100110101011;
		16'b0000110000111001 : data_out =  24'b000000000100100110111110;
		16'b0000110000111011 : data_out =  24'b000000000100100111010001;
		16'b0000110000111101 : data_out =  24'b000000000100100111100100;
		16'b0000110000111111 : data_out =  24'b000000000100100111110110;
		16'b0000110001000001 : data_out =  24'b000000000100101000001001;
		16'b0000110001000011 : data_out =  24'b000000000100101000011100;
		16'b0000110001000101 : data_out =  24'b000000000100101000101111;
		16'b0000110001000111 : data_out =  24'b000000000100101001000010;
		16'b0000110001001001 : data_out =  24'b000000000100101001010101;
		16'b0000110001001011 : data_out =  24'b000000000100101001101000;
		16'b0000110001001101 : data_out =  24'b000000000100101001111011;
		16'b0000110001001111 : data_out =  24'b000000000100101010001111;
		16'b0000110001010001 : data_out =  24'b000000000100101010100010;
		16'b0000110001010011 : data_out =  24'b000000000100101010110101;
		16'b0000110001010110 : data_out =  24'b000000000100101011001000;
		16'b0000110001011000 : data_out =  24'b000000000100101011011011;
		16'b0000110001011010 : data_out =  24'b000000000100101011101110;
		16'b0000110001011100 : data_out =  24'b000000000100101100000001;
		16'b0000110001011110 : data_out =  24'b000000000100101100010101;
		16'b0000110001100000 : data_out =  24'b000000000100101100101000;
		16'b0000110001100010 : data_out =  24'b000000000100101100111011;
		16'b0000110001100100 : data_out =  24'b000000000100101101001110;
		16'b0000110001100110 : data_out =  24'b000000000100101101100010;
		16'b0000110001101000 : data_out =  24'b000000000100101101110101;
		16'b0000110001101010 : data_out =  24'b000000000100101110001000;
		16'b0000110001101100 : data_out =  24'b000000000100101110011100;
		16'b0000110001101110 : data_out =  24'b000000000100101110101111;
		16'b0000110001110000 : data_out =  24'b000000000100101111000010;
		16'b0000110001110010 : data_out =  24'b000000000100101111010110;
		16'b0000110001110100 : data_out =  24'b000000000100101111101001;
		16'b0000110001110110 : data_out =  24'b000000000100101111111101;
		16'b0000110001111000 : data_out =  24'b000000000100110000010000;
		16'b0000110001111010 : data_out =  24'b000000000100110000100100;
		16'b0000110001111100 : data_out =  24'b000000000100110000110111;
		16'b0000110001111110 : data_out =  24'b000000000100110001001011;
		16'b0000110010000001 : data_out =  24'b000000000100110001011110;
		16'b0000110010000011 : data_out =  24'b000000000100110001110010;
		16'b0000110010000101 : data_out =  24'b000000000100110010000101;
		16'b0000110010000111 : data_out =  24'b000000000100110010011001;
		16'b0000110010001001 : data_out =  24'b000000000100110010101101;
		16'b0000110010001011 : data_out =  24'b000000000100110011000000;
		16'b0000110010001101 : data_out =  24'b000000000100110011010100;
		16'b0000110010001111 : data_out =  24'b000000000100110011101000;
		16'b0000110010010001 : data_out =  24'b000000000100110011111011;
		16'b0000110010010011 : data_out =  24'b000000000100110100001111;
		16'b0000110010010101 : data_out =  24'b000000000100110100100011;
		16'b0000110010010111 : data_out =  24'b000000000100110100110110;
		16'b0000110010011001 : data_out =  24'b000000000100110101001010;
		16'b0000110010011011 : data_out =  24'b000000000100110101011110;
		16'b0000110010011101 : data_out =  24'b000000000100110101110010;
		16'b0000110010011111 : data_out =  24'b000000000100110110000110;
		16'b0000110010100001 : data_out =  24'b000000000100110110011010;
		16'b0000110010100011 : data_out =  24'b000000000100110110101101;
		16'b0000110010100101 : data_out =  24'b000000000100110111000001;
		16'b0000110010100111 : data_out =  24'b000000000100110111010101;
		16'b0000110010101001 : data_out =  24'b000000000100110111101001;
		16'b0000110010101100 : data_out =  24'b000000000100110111111101;
		16'b0000110010101110 : data_out =  24'b000000000100111000010001;
		16'b0000110010110000 : data_out =  24'b000000000100111000100101;
		16'b0000110010110010 : data_out =  24'b000000000100111000111001;
		16'b0000110010110100 : data_out =  24'b000000000100111001001101;
		16'b0000110010110110 : data_out =  24'b000000000100111001100001;
		16'b0000110010111000 : data_out =  24'b000000000100111001110101;
		16'b0000110010111010 : data_out =  24'b000000000100111010001001;
		16'b0000110010111100 : data_out =  24'b000000000100111010011101;
		16'b0000110010111110 : data_out =  24'b000000000100111010110010;
		16'b0000110011000000 : data_out =  24'b000000000100111011000110;
		16'b0000110011000010 : data_out =  24'b000000000100111011011010;
		16'b0000110011000100 : data_out =  24'b000000000100111011101110;
		16'b0000110011000110 : data_out =  24'b000000000100111100000010;
		16'b0000110011001000 : data_out =  24'b000000000100111100010111;
		16'b0000110011001010 : data_out =  24'b000000000100111100101011;
		16'b0000110011001100 : data_out =  24'b000000000100111100111111;
		16'b0000110011001110 : data_out =  24'b000000000100111101010011;
		16'b0000110011010000 : data_out =  24'b000000000100111101101000;
		16'b0000110011010010 : data_out =  24'b000000000100111101111100;
		16'b0000110011010100 : data_out =  24'b000000000100111110010000;
		16'b0000110011010111 : data_out =  24'b000000000100111110100101;
		16'b0000110011011001 : data_out =  24'b000000000100111110111001;
		16'b0000110011011011 : data_out =  24'b000000000100111111001110;
		16'b0000110011011101 : data_out =  24'b000000000100111111100010;
		16'b0000110011011111 : data_out =  24'b000000000100111111110111;
		16'b0000110011100001 : data_out =  24'b000000000101000000001011;
		16'b0000110011100011 : data_out =  24'b000000000101000000100000;
		16'b0000110011100101 : data_out =  24'b000000000101000000110100;
		16'b0000110011100111 : data_out =  24'b000000000101000001001001;
		16'b0000110011101001 : data_out =  24'b000000000101000001011101;
		16'b0000110011101011 : data_out =  24'b000000000101000001110010;
		16'b0000110011101101 : data_out =  24'b000000000101000010000110;
		16'b0000110011101111 : data_out =  24'b000000000101000010011011;
		16'b0000110011110001 : data_out =  24'b000000000101000010110000;
		16'b0000110011110011 : data_out =  24'b000000000101000011000100;
		16'b0000110011110101 : data_out =  24'b000000000101000011011001;
		16'b0000110011110111 : data_out =  24'b000000000101000011101110;
		16'b0000110011111001 : data_out =  24'b000000000101000100000010;
		16'b0000110011111011 : data_out =  24'b000000000101000100010111;
		16'b0000110011111101 : data_out =  24'b000000000101000100101100;
		16'b0000110011111111 : data_out =  24'b000000000101000101000001;
		16'b0000110100000010 : data_out =  24'b000000000101000101010110;
		16'b0000110100000100 : data_out =  24'b000000000101000101101010;
		16'b0000110100000110 : data_out =  24'b000000000101000101111111;
		16'b0000110100001000 : data_out =  24'b000000000101000110010100;
		16'b0000110100001010 : data_out =  24'b000000000101000110101001;
		16'b0000110100001100 : data_out =  24'b000000000101000110111110;
		16'b0000110100001110 : data_out =  24'b000000000101000111010011;
		16'b0000110100010000 : data_out =  24'b000000000101000111101000;
		16'b0000110100010010 : data_out =  24'b000000000101000111111101;
		16'b0000110100010100 : data_out =  24'b000000000101001000010010;
		16'b0000110100010110 : data_out =  24'b000000000101001000100111;
		16'b0000110100011000 : data_out =  24'b000000000101001000111100;
		16'b0000110100011010 : data_out =  24'b000000000101001001010001;
		16'b0000110100011100 : data_out =  24'b000000000101001001100110;
		16'b0000110100011110 : data_out =  24'b000000000101001001111011;
		16'b0000110100100000 : data_out =  24'b000000000101001010010000;
		16'b0000110100100010 : data_out =  24'b000000000101001010100101;
		16'b0000110100100100 : data_out =  24'b000000000101001010111011;
		16'b0000110100100110 : data_out =  24'b000000000101001011010000;
		16'b0000110100101000 : data_out =  24'b000000000101001011100101;
		16'b0000110100101011 : data_out =  24'b000000000101001011111010;
		16'b0000110100101101 : data_out =  24'b000000000101001100001111;
		16'b0000110100101111 : data_out =  24'b000000000101001100100101;
		16'b0000110100110001 : data_out =  24'b000000000101001100111010;
		16'b0000110100110011 : data_out =  24'b000000000101001101001111;
		16'b0000110100110101 : data_out =  24'b000000000101001101100101;
		16'b0000110100110111 : data_out =  24'b000000000101001101111010;
		16'b0000110100111001 : data_out =  24'b000000000101001110001111;
		16'b0000110100111011 : data_out =  24'b000000000101001110100101;
		16'b0000110100111101 : data_out =  24'b000000000101001110111010;
		16'b0000110100111111 : data_out =  24'b000000000101001111010000;
		16'b0000110101000001 : data_out =  24'b000000000101001111100101;
		16'b0000110101000011 : data_out =  24'b000000000101001111111011;
		16'b0000110101000101 : data_out =  24'b000000000101010000010000;
		16'b0000110101000111 : data_out =  24'b000000000101010000100110;
		16'b0000110101001001 : data_out =  24'b000000000101010000111011;
		16'b0000110101001011 : data_out =  24'b000000000101010001010001;
		16'b0000110101001101 : data_out =  24'b000000000101010001100110;
		16'b0000110101001111 : data_out =  24'b000000000101010001111100;
		16'b0000110101010001 : data_out =  24'b000000000101010010010010;
		16'b0000110101010011 : data_out =  24'b000000000101010010100111;
		16'b0000110101010110 : data_out =  24'b000000000101010010111101;
		16'b0000110101011000 : data_out =  24'b000000000101010011010011;
		16'b0000110101011010 : data_out =  24'b000000000101010011101000;
		16'b0000110101011100 : data_out =  24'b000000000101010011111110;
		16'b0000110101011110 : data_out =  24'b000000000101010100010100;
		16'b0000110101100000 : data_out =  24'b000000000101010100101010;
		16'b0000110101100010 : data_out =  24'b000000000101010101000000;
		16'b0000110101100100 : data_out =  24'b000000000101010101010101;
		16'b0000110101100110 : data_out =  24'b000000000101010101101011;
		16'b0000110101101000 : data_out =  24'b000000000101010110000001;
		16'b0000110101101010 : data_out =  24'b000000000101010110010111;
		16'b0000110101101100 : data_out =  24'b000000000101010110101101;
		16'b0000110101101110 : data_out =  24'b000000000101010111000011;
		16'b0000110101110000 : data_out =  24'b000000000101010111011001;
		16'b0000110101110010 : data_out =  24'b000000000101010111101111;
		16'b0000110101110100 : data_out =  24'b000000000101011000000101;
		16'b0000110101110110 : data_out =  24'b000000000101011000011011;
		16'b0000110101111000 : data_out =  24'b000000000101011000110001;
		16'b0000110101111010 : data_out =  24'b000000000101011001000111;
		16'b0000110101111100 : data_out =  24'b000000000101011001011101;
		16'b0000110101111110 : data_out =  24'b000000000101011001110011;
		16'b0000110110000001 : data_out =  24'b000000000101011010001001;
		16'b0000110110000011 : data_out =  24'b000000000101011010100000;
		16'b0000110110000101 : data_out =  24'b000000000101011010110110;
		16'b0000110110000111 : data_out =  24'b000000000101011011001100;
		16'b0000110110001001 : data_out =  24'b000000000101011011100010;
		16'b0000110110001011 : data_out =  24'b000000000101011011111000;
		16'b0000110110001101 : data_out =  24'b000000000101011100001111;
		16'b0000110110001111 : data_out =  24'b000000000101011100100101;
		16'b0000110110010001 : data_out =  24'b000000000101011100111011;
		16'b0000110110010011 : data_out =  24'b000000000101011101010010;
		16'b0000110110010101 : data_out =  24'b000000000101011101101000;
		16'b0000110110010111 : data_out =  24'b000000000101011101111110;
		16'b0000110110011001 : data_out =  24'b000000000101011110010101;
		16'b0000110110011011 : data_out =  24'b000000000101011110101011;
		16'b0000110110011101 : data_out =  24'b000000000101011111000010;
		16'b0000110110011111 : data_out =  24'b000000000101011111011000;
		16'b0000110110100001 : data_out =  24'b000000000101011111101111;
		16'b0000110110100011 : data_out =  24'b000000000101100000000101;
		16'b0000110110100101 : data_out =  24'b000000000101100000011100;
		16'b0000110110100111 : data_out =  24'b000000000101100000110010;
		16'b0000110110101001 : data_out =  24'b000000000101100001001001;
		16'b0000110110101100 : data_out =  24'b000000000101100001011111;
		16'b0000110110101110 : data_out =  24'b000000000101100001110110;
		16'b0000110110110000 : data_out =  24'b000000000101100010001101;
		16'b0000110110110010 : data_out =  24'b000000000101100010100011;
		16'b0000110110110100 : data_out =  24'b000000000101100010111010;
		16'b0000110110110110 : data_out =  24'b000000000101100011010001;
		16'b0000110110111000 : data_out =  24'b000000000101100011101000;
		16'b0000110110111010 : data_out =  24'b000000000101100011111110;
		16'b0000110110111100 : data_out =  24'b000000000101100100010101;
		16'b0000110110111110 : data_out =  24'b000000000101100100101100;
		16'b0000110111000000 : data_out =  24'b000000000101100101000011;
		16'b0000110111000010 : data_out =  24'b000000000101100101011010;
		16'b0000110111000100 : data_out =  24'b000000000101100101110001;
		16'b0000110111000110 : data_out =  24'b000000000101100110001000;
		16'b0000110111001000 : data_out =  24'b000000000101100110011110;
		16'b0000110111001010 : data_out =  24'b000000000101100110110101;
		16'b0000110111001100 : data_out =  24'b000000000101100111001100;
		16'b0000110111001110 : data_out =  24'b000000000101100111100011;
		16'b0000110111010000 : data_out =  24'b000000000101100111111010;
		16'b0000110111010010 : data_out =  24'b000000000101101000010001;
		16'b0000110111010100 : data_out =  24'b000000000101101000101001;
		16'b0000110111010111 : data_out =  24'b000000000101101001000000;
		16'b0000110111011001 : data_out =  24'b000000000101101001010111;
		16'b0000110111011011 : data_out =  24'b000000000101101001101110;
		16'b0000110111011101 : data_out =  24'b000000000101101010000101;
		16'b0000110111011111 : data_out =  24'b000000000101101010011100;
		16'b0000110111100001 : data_out =  24'b000000000101101010110011;
		16'b0000110111100011 : data_out =  24'b000000000101101011001011;
		16'b0000110111100101 : data_out =  24'b000000000101101011100010;
		16'b0000110111100111 : data_out =  24'b000000000101101011111001;
		16'b0000110111101001 : data_out =  24'b000000000101101100010000;
		16'b0000110111101011 : data_out =  24'b000000000101101100101000;
		16'b0000110111101101 : data_out =  24'b000000000101101100111111;
		16'b0000110111101111 : data_out =  24'b000000000101101101010111;
		16'b0000110111110001 : data_out =  24'b000000000101101101101110;
		16'b0000110111110011 : data_out =  24'b000000000101101110000101;
		16'b0000110111110101 : data_out =  24'b000000000101101110011101;
		16'b0000110111110111 : data_out =  24'b000000000101101110110100;
		16'b0000110111111001 : data_out =  24'b000000000101101111001100;
		16'b0000110111111011 : data_out =  24'b000000000101101111100011;
		16'b0000110111111101 : data_out =  24'b000000000101101111111011;
		16'b0000110111111111 : data_out =  24'b000000000101110000010010;
		16'b0000111000000010 : data_out =  24'b000000000101110000101010;
		16'b0000111000000100 : data_out =  24'b000000000101110001000010;
		16'b0000111000000110 : data_out =  24'b000000000101110001011001;
		16'b0000111000001000 : data_out =  24'b000000000101110001110001;
		16'b0000111000001010 : data_out =  24'b000000000101110010001001;
		16'b0000111000001100 : data_out =  24'b000000000101110010100000;
		16'b0000111000001110 : data_out =  24'b000000000101110010111000;
		16'b0000111000010000 : data_out =  24'b000000000101110011010000;
		16'b0000111000010010 : data_out =  24'b000000000101110011100111;
		16'b0000111000010100 : data_out =  24'b000000000101110011111111;
		16'b0000111000010110 : data_out =  24'b000000000101110100010111;
		16'b0000111000011000 : data_out =  24'b000000000101110100101111;
		16'b0000111000011010 : data_out =  24'b000000000101110101000111;
		16'b0000111000011100 : data_out =  24'b000000000101110101011111;
		16'b0000111000011110 : data_out =  24'b000000000101110101110111;
		16'b0000111000100000 : data_out =  24'b000000000101110110001111;
		16'b0000111000100010 : data_out =  24'b000000000101110110100110;
		16'b0000111000100100 : data_out =  24'b000000000101110110111110;
		16'b0000111000100110 : data_out =  24'b000000000101110111010110;
		16'b0000111000101000 : data_out =  24'b000000000101110111101111;
		16'b0000111000101011 : data_out =  24'b000000000101111000000111;
		16'b0000111000101101 : data_out =  24'b000000000101111000011111;
		16'b0000111000101111 : data_out =  24'b000000000101111000110111;
		16'b0000111000110001 : data_out =  24'b000000000101111001001111;
		16'b0000111000110011 : data_out =  24'b000000000101111001100111;
		16'b0000111000110101 : data_out =  24'b000000000101111001111111;
		16'b0000111000110111 : data_out =  24'b000000000101111010010111;
		16'b0000111000111001 : data_out =  24'b000000000101111010110000;
		16'b0000111000111011 : data_out =  24'b000000000101111011001000;
		16'b0000111000111101 : data_out =  24'b000000000101111011100000;
		16'b0000111000111111 : data_out =  24'b000000000101111011111000;
		16'b0000111001000001 : data_out =  24'b000000000101111100010001;
		16'b0000111001000011 : data_out =  24'b000000000101111100101001;
		16'b0000111001000101 : data_out =  24'b000000000101111101000010;
		16'b0000111001000111 : data_out =  24'b000000000101111101011010;
		16'b0000111001001001 : data_out =  24'b000000000101111101110010;
		16'b0000111001001011 : data_out =  24'b000000000101111110001011;
		16'b0000111001001101 : data_out =  24'b000000000101111110100011;
		16'b0000111001001111 : data_out =  24'b000000000101111110111100;
		16'b0000111001010001 : data_out =  24'b000000000101111111010100;
		16'b0000111001010011 : data_out =  24'b000000000101111111101101;
		16'b0000111001010110 : data_out =  24'b000000000110000000000101;
		16'b0000111001011000 : data_out =  24'b000000000110000000011110;
		16'b0000111001011010 : data_out =  24'b000000000110000000110111;
		16'b0000111001011100 : data_out =  24'b000000000110000001001111;
		16'b0000111001011110 : data_out =  24'b000000000110000001101000;
		16'b0000111001100000 : data_out =  24'b000000000110000010000001;
		16'b0000111001100010 : data_out =  24'b000000000110000010011001;
		16'b0000111001100100 : data_out =  24'b000000000110000010110010;
		16'b0000111001100110 : data_out =  24'b000000000110000011001011;
		16'b0000111001101000 : data_out =  24'b000000000110000011100100;
		16'b0000111001101010 : data_out =  24'b000000000110000011111100;
		16'b0000111001101100 : data_out =  24'b000000000110000100010101;
		16'b0000111001101110 : data_out =  24'b000000000110000100101110;
		16'b0000111001110000 : data_out =  24'b000000000110000101000111;
		16'b0000111001110010 : data_out =  24'b000000000110000101100000;
		16'b0000111001110100 : data_out =  24'b000000000110000101111001;
		16'b0000111001110110 : data_out =  24'b000000000110000110010010;
		16'b0000111001111000 : data_out =  24'b000000000110000110101011;
		16'b0000111001111010 : data_out =  24'b000000000110000111000100;
		16'b0000111001111100 : data_out =  24'b000000000110000111011101;
		16'b0000111001111110 : data_out =  24'b000000000110000111110110;
		16'b0000111010000001 : data_out =  24'b000000000110001000001111;
		16'b0000111010000011 : data_out =  24'b000000000110001000101000;
		16'b0000111010000101 : data_out =  24'b000000000110001001000001;
		16'b0000111010000111 : data_out =  24'b000000000110001001011011;
		16'b0000111010001001 : data_out =  24'b000000000110001001110100;
		16'b0000111010001011 : data_out =  24'b000000000110001010001101;
		16'b0000111010001101 : data_out =  24'b000000000110001010100110;
		16'b0000111010001111 : data_out =  24'b000000000110001010111111;
		16'b0000111010010001 : data_out =  24'b000000000110001011011001;
		16'b0000111010010011 : data_out =  24'b000000000110001011110010;
		16'b0000111010010101 : data_out =  24'b000000000110001100001011;
		16'b0000111010010111 : data_out =  24'b000000000110001100100101;
		16'b0000111010011001 : data_out =  24'b000000000110001100111110;
		16'b0000111010011011 : data_out =  24'b000000000110001101011000;
		16'b0000111010011101 : data_out =  24'b000000000110001101110001;
		16'b0000111010011111 : data_out =  24'b000000000110001110001010;
		16'b0000111010100001 : data_out =  24'b000000000110001110100100;
		16'b0000111010100011 : data_out =  24'b000000000110001110111101;
		16'b0000111010100101 : data_out =  24'b000000000110001111010111;
		16'b0000111010100111 : data_out =  24'b000000000110001111110001;
		16'b0000111010101001 : data_out =  24'b000000000110010000001010;
		16'b0000111010101100 : data_out =  24'b000000000110010000100100;
		16'b0000111010101110 : data_out =  24'b000000000110010000111101;
		16'b0000111010110000 : data_out =  24'b000000000110010001010111;
		16'b0000111010110010 : data_out =  24'b000000000110010001110001;
		16'b0000111010110100 : data_out =  24'b000000000110010010001011;
		16'b0000111010110110 : data_out =  24'b000000000110010010100100;
		16'b0000111010111000 : data_out =  24'b000000000110010010111110;
		16'b0000111010111010 : data_out =  24'b000000000110010011011000;
		16'b0000111010111100 : data_out =  24'b000000000110010011110010;
		16'b0000111010111110 : data_out =  24'b000000000110010100001100;
		16'b0000111011000000 : data_out =  24'b000000000110010100100101;
		16'b0000111011000010 : data_out =  24'b000000000110010100111111;
		16'b0000111011000100 : data_out =  24'b000000000110010101011001;
		16'b0000111011000110 : data_out =  24'b000000000110010101110011;
		16'b0000111011001000 : data_out =  24'b000000000110010110001101;
		16'b0000111011001010 : data_out =  24'b000000000110010110100111;
		16'b0000111011001100 : data_out =  24'b000000000110010111000001;
		16'b0000111011001110 : data_out =  24'b000000000110010111011011;
		16'b0000111011010000 : data_out =  24'b000000000110010111110101;
		16'b0000111011010010 : data_out =  24'b000000000110011000010000;
		16'b0000111011010100 : data_out =  24'b000000000110011000101010;
		16'b0000111011010111 : data_out =  24'b000000000110011001000100;
		16'b0000111011011001 : data_out =  24'b000000000110011001011110;
		16'b0000111011011011 : data_out =  24'b000000000110011001111000;
		16'b0000111011011101 : data_out =  24'b000000000110011010010011;
		16'b0000111011011111 : data_out =  24'b000000000110011010101101;
		16'b0000111011100001 : data_out =  24'b000000000110011011000111;
		16'b0000111011100011 : data_out =  24'b000000000110011011100001;
		16'b0000111011100101 : data_out =  24'b000000000110011011111100;
		16'b0000111011100111 : data_out =  24'b000000000110011100010110;
		16'b0000111011101001 : data_out =  24'b000000000110011100110001;
		16'b0000111011101011 : data_out =  24'b000000000110011101001011;
		16'b0000111011101101 : data_out =  24'b000000000110011101100101;
		16'b0000111011101111 : data_out =  24'b000000000110011110000000;
		16'b0000111011110001 : data_out =  24'b000000000110011110011010;
		16'b0000111011110011 : data_out =  24'b000000000110011110110101;
		16'b0000111011110101 : data_out =  24'b000000000110011111010000;
		16'b0000111011110111 : data_out =  24'b000000000110011111101010;
		16'b0000111011111001 : data_out =  24'b000000000110100000000101;
		16'b0000111011111011 : data_out =  24'b000000000110100000011111;
		16'b0000111011111101 : data_out =  24'b000000000110100000111010;
		16'b0000111011111111 : data_out =  24'b000000000110100001010101;
		16'b0000111100000010 : data_out =  24'b000000000110100001101111;
		16'b0000111100000100 : data_out =  24'b000000000110100010001010;
		16'b0000111100000110 : data_out =  24'b000000000110100010100101;
		16'b0000111100001000 : data_out =  24'b000000000110100011000000;
		16'b0000111100001010 : data_out =  24'b000000000110100011011011;
		16'b0000111100001100 : data_out =  24'b000000000110100011110110;
		16'b0000111100001110 : data_out =  24'b000000000110100100010000;
		16'b0000111100010000 : data_out =  24'b000000000110100100101011;
		16'b0000111100010010 : data_out =  24'b000000000110100101000110;
		16'b0000111100010100 : data_out =  24'b000000000110100101100001;
		16'b0000111100010110 : data_out =  24'b000000000110100101111100;
		16'b0000111100011000 : data_out =  24'b000000000110100110010111;
		16'b0000111100011010 : data_out =  24'b000000000110100110110010;
		16'b0000111100011100 : data_out =  24'b000000000110100111001101;
		16'b0000111100011110 : data_out =  24'b000000000110100111101000;
		16'b0000111100100000 : data_out =  24'b000000000110101000000100;
		16'b0000111100100010 : data_out =  24'b000000000110101000011111;
		16'b0000111100100100 : data_out =  24'b000000000110101000111010;
		16'b0000111100100110 : data_out =  24'b000000000110101001010101;
		16'b0000111100101000 : data_out =  24'b000000000110101001110000;
		16'b0000111100101011 : data_out =  24'b000000000110101010001100;
		16'b0000111100101101 : data_out =  24'b000000000110101010100111;
		16'b0000111100101111 : data_out =  24'b000000000110101011000010;
		16'b0000111100110001 : data_out =  24'b000000000110101011011110;
		16'b0000111100110011 : data_out =  24'b000000000110101011111001;
		16'b0000111100110101 : data_out =  24'b000000000110101100010100;
		16'b0000111100110111 : data_out =  24'b000000000110101100110000;
		16'b0000111100111001 : data_out =  24'b000000000110101101001011;
		16'b0000111100111011 : data_out =  24'b000000000110101101100111;
		16'b0000111100111101 : data_out =  24'b000000000110101110000010;
		16'b0000111100111111 : data_out =  24'b000000000110101110011110;
		16'b0000111101000001 : data_out =  24'b000000000110101110111001;
		16'b0000111101000011 : data_out =  24'b000000000110101111010101;
		16'b0000111101000101 : data_out =  24'b000000000110101111110001;
		16'b0000111101000111 : data_out =  24'b000000000110110000001100;
		16'b0000111101001001 : data_out =  24'b000000000110110000101000;
		16'b0000111101001011 : data_out =  24'b000000000110110001000100;
		16'b0000111101001101 : data_out =  24'b000000000110110001011111;
		16'b0000111101001111 : data_out =  24'b000000000110110001111011;
		16'b0000111101010001 : data_out =  24'b000000000110110010010111;
		16'b0000111101010011 : data_out =  24'b000000000110110010110011;
		16'b0000111101010110 : data_out =  24'b000000000110110011001110;
		16'b0000111101011000 : data_out =  24'b000000000110110011101010;
		16'b0000111101011010 : data_out =  24'b000000000110110100000110;
		16'b0000111101011100 : data_out =  24'b000000000110110100100010;
		16'b0000111101011110 : data_out =  24'b000000000110110100111110;
		16'b0000111101100000 : data_out =  24'b000000000110110101011010;
		16'b0000111101100010 : data_out =  24'b000000000110110101110110;
		16'b0000111101100100 : data_out =  24'b000000000110110110010010;
		16'b0000111101100110 : data_out =  24'b000000000110110110101110;
		16'b0000111101101000 : data_out =  24'b000000000110110111001010;
		16'b0000111101101010 : data_out =  24'b000000000110110111100110;
		16'b0000111101101100 : data_out =  24'b000000000110111000000011;
		16'b0000111101101110 : data_out =  24'b000000000110111000011111;
		16'b0000111101110000 : data_out =  24'b000000000110111000111011;
		16'b0000111101110010 : data_out =  24'b000000000110111001010111;
		16'b0000111101110100 : data_out =  24'b000000000110111001110011;
		16'b0000111101110110 : data_out =  24'b000000000110111010010000;
		16'b0000111101111000 : data_out =  24'b000000000110111010101100;
		16'b0000111101111010 : data_out =  24'b000000000110111011001000;
		16'b0000111101111100 : data_out =  24'b000000000110111011100101;
		16'b0000111101111110 : data_out =  24'b000000000110111100000001;
		16'b0000111110000001 : data_out =  24'b000000000110111100011110;
		16'b0000111110000011 : data_out =  24'b000000000110111100111010;
		16'b0000111110000101 : data_out =  24'b000000000110111101010111;
		16'b0000111110000111 : data_out =  24'b000000000110111101110011;
		16'b0000111110001001 : data_out =  24'b000000000110111110010000;
		16'b0000111110001011 : data_out =  24'b000000000110111110101100;
		16'b0000111110001101 : data_out =  24'b000000000110111111001001;
		16'b0000111110001111 : data_out =  24'b000000000110111111100101;
		16'b0000111110010001 : data_out =  24'b000000000111000000000010;
		16'b0000111110010011 : data_out =  24'b000000000111000000011111;
		16'b0000111110010101 : data_out =  24'b000000000111000000111011;
		16'b0000111110010111 : data_out =  24'b000000000111000001011000;
		16'b0000111110011001 : data_out =  24'b000000000111000001110101;
		16'b0000111110011011 : data_out =  24'b000000000111000010010010;
		16'b0000111110011101 : data_out =  24'b000000000111000010101111;
		16'b0000111110011111 : data_out =  24'b000000000111000011001100;
		16'b0000111110100001 : data_out =  24'b000000000111000011101000;
		16'b0000111110100011 : data_out =  24'b000000000111000100000101;
		16'b0000111110100101 : data_out =  24'b000000000111000100100010;
		16'b0000111110100111 : data_out =  24'b000000000111000100111111;
		16'b0000111110101001 : data_out =  24'b000000000111000101011100;
		16'b0000111110101100 : data_out =  24'b000000000111000101111001;
		16'b0000111110101110 : data_out =  24'b000000000111000110010110;
		16'b0000111110110000 : data_out =  24'b000000000111000110110011;
		16'b0000111110110010 : data_out =  24'b000000000111000111010001;
		16'b0000111110110100 : data_out =  24'b000000000111000111101110;
		16'b0000111110110110 : data_out =  24'b000000000111001000001011;
		16'b0000111110111000 : data_out =  24'b000000000111001000101000;
		16'b0000111110111010 : data_out =  24'b000000000111001001000101;
		16'b0000111110111100 : data_out =  24'b000000000111001001100011;
		16'b0000111110111110 : data_out =  24'b000000000111001010000000;
		16'b0000111111000000 : data_out =  24'b000000000111001010011101;
		16'b0000111111000010 : data_out =  24'b000000000111001010111011;
		16'b0000111111000100 : data_out =  24'b000000000111001011011000;
		16'b0000111111000110 : data_out =  24'b000000000111001011110101;
		16'b0000111111001000 : data_out =  24'b000000000111001100010011;
		16'b0000111111001010 : data_out =  24'b000000000111001100110000;
		16'b0000111111001100 : data_out =  24'b000000000111001101001110;
		16'b0000111111001110 : data_out =  24'b000000000111001101101011;
		16'b0000111111010000 : data_out =  24'b000000000111001110001001;
		16'b0000111111010010 : data_out =  24'b000000000111001110100111;
		16'b0000111111010100 : data_out =  24'b000000000111001111000100;
		16'b0000111111010111 : data_out =  24'b000000000111001111100010;
		16'b0000111111011001 : data_out =  24'b000000000111001111111111;
		16'b0000111111011011 : data_out =  24'b000000000111010000011101;
		16'b0000111111011101 : data_out =  24'b000000000111010000111011;
		16'b0000111111011111 : data_out =  24'b000000000111010001011001;
		16'b0000111111100001 : data_out =  24'b000000000111010001110110;
		16'b0000111111100011 : data_out =  24'b000000000111010010010100;
		16'b0000111111100101 : data_out =  24'b000000000111010010110010;
		16'b0000111111100111 : data_out =  24'b000000000111010011010000;
		16'b0000111111101001 : data_out =  24'b000000000111010011101110;
		16'b0000111111101011 : data_out =  24'b000000000111010100001100;
		16'b0000111111101101 : data_out =  24'b000000000111010100101010;
		16'b0000111111101111 : data_out =  24'b000000000111010101001000;
		16'b0000111111110001 : data_out =  24'b000000000111010101100110;
		16'b0000111111110011 : data_out =  24'b000000000111010110000100;
		16'b0000111111110101 : data_out =  24'b000000000111010110100010;
		16'b0000111111110111 : data_out =  24'b000000000111010111000000;
		16'b0000111111111001 : data_out =  24'b000000000111010111011110;
		16'b0000111111111011 : data_out =  24'b000000000111010111111101;
		16'b0000111111111101 : data_out =  24'b000000000111011000011011;
		16'b0000111111111111 : data_out =  24'b000000000111011000111001;
		16'b0001000000000010 : data_out =  24'b000000000111011001010111;
		16'b0001000000000100 : data_out =  24'b000000000111011001110110;
		16'b0001000000000110 : data_out =  24'b000000000111011010010100;
		16'b0001000000001000 : data_out =  24'b000000000111011010110010;
		16'b0001000000001010 : data_out =  24'b000000000111011011010001;
		16'b0001000000001100 : data_out =  24'b000000000111011011101111;
		16'b0001000000001110 : data_out =  24'b000000000111011100001110;
		16'b0001000000010000 : data_out =  24'b000000000111011100101100;
		16'b0001000000010010 : data_out =  24'b000000000111011101001011;
		16'b0001000000010100 : data_out =  24'b000000000111011101101001;
		16'b0001000000010110 : data_out =  24'b000000000111011110001000;
		16'b0001000000011000 : data_out =  24'b000000000111011110100110;
		16'b0001000000011010 : data_out =  24'b000000000111011111000101;
		16'b0001000000011100 : data_out =  24'b000000000111011111100100;
		16'b0001000000011110 : data_out =  24'b000000000111100000000010;
		16'b0001000000100000 : data_out =  24'b000000000111100000100001;
		16'b0001000000100010 : data_out =  24'b000000000111100001000000;
		16'b0001000000100100 : data_out =  24'b000000000111100001011111;
		16'b0001000000100110 : data_out =  24'b000000000111100001111110;
		16'b0001000000101000 : data_out =  24'b000000000111100010011100;
		16'b0001000000101011 : data_out =  24'b000000000111100010111011;
		16'b0001000000101101 : data_out =  24'b000000000111100011011010;
		16'b0001000000101111 : data_out =  24'b000000000111100011111001;
		16'b0001000000110001 : data_out =  24'b000000000111100100011000;
		16'b0001000000110011 : data_out =  24'b000000000111100100110111;
		16'b0001000000110101 : data_out =  24'b000000000111100101010110;
		16'b0001000000110111 : data_out =  24'b000000000111100101110101;
		16'b0001000000111001 : data_out =  24'b000000000111100110010100;
		16'b0001000000111011 : data_out =  24'b000000000111100110110100;
		16'b0001000000111101 : data_out =  24'b000000000111100111010011;
		16'b0001000000111111 : data_out =  24'b000000000111100111110010;
		16'b0001000001000001 : data_out =  24'b000000000111101000010001;
		16'b0001000001000011 : data_out =  24'b000000000111101000110001;
		16'b0001000001000101 : data_out =  24'b000000000111101001010000;
		16'b0001000001000111 : data_out =  24'b000000000111101001101111;
		16'b0001000001001001 : data_out =  24'b000000000111101010001110;
		16'b0001000001001011 : data_out =  24'b000000000111101010101110;
		16'b0001000001001101 : data_out =  24'b000000000111101011001101;
		16'b0001000001001111 : data_out =  24'b000000000111101011101101;
		16'b0001000001010001 : data_out =  24'b000000000111101100001100;
		16'b0001000001010011 : data_out =  24'b000000000111101100101100;
		16'b0001000001010110 : data_out =  24'b000000000111101101001011;
		16'b0001000001011000 : data_out =  24'b000000000111101101101011;
		16'b0001000001011010 : data_out =  24'b000000000111101110001010;
		16'b0001000001011100 : data_out =  24'b000000000111101110101010;
		16'b0001000001011110 : data_out =  24'b000000000111101111001010;
		16'b0001000001100000 : data_out =  24'b000000000111101111101010;
		16'b0001000001100010 : data_out =  24'b000000000111110000001001;
		16'b0001000001100100 : data_out =  24'b000000000111110000101001;
		16'b0001000001100110 : data_out =  24'b000000000111110001001001;
		16'b0001000001101000 : data_out =  24'b000000000111110001101001;
		16'b0001000001101010 : data_out =  24'b000000000111110010001001;
		16'b0001000001101100 : data_out =  24'b000000000111110010101000;
		16'b0001000001101110 : data_out =  24'b000000000111110011001000;
		16'b0001000001110000 : data_out =  24'b000000000111110011101000;
		16'b0001000001110010 : data_out =  24'b000000000111110100001000;
		16'b0001000001110100 : data_out =  24'b000000000111110100101000;
		16'b0001000001110110 : data_out =  24'b000000000111110101001000;
		16'b0001000001111000 : data_out =  24'b000000000111110101101000;
		16'b0001000001111010 : data_out =  24'b000000000111110110001001;
		16'b0001000001111100 : data_out =  24'b000000000111110110101001;
		16'b0001000001111110 : data_out =  24'b000000000111110111001001;
		16'b0001000010000001 : data_out =  24'b000000000111110111101001;
		16'b0001000010000011 : data_out =  24'b000000000111111000001001;
		16'b0001000010000101 : data_out =  24'b000000000111111000101010;
		16'b0001000010000111 : data_out =  24'b000000000111111001001010;
		16'b0001000010001001 : data_out =  24'b000000000111111001101010;
		16'b0001000010001011 : data_out =  24'b000000000111111010001011;
		16'b0001000010001101 : data_out =  24'b000000000111111010101011;
		16'b0001000010001111 : data_out =  24'b000000000111111011001100;
		16'b0001000010010001 : data_out =  24'b000000000111111011101100;
		16'b0001000010010011 : data_out =  24'b000000000111111100001101;
		16'b0001000010010101 : data_out =  24'b000000000111111100101101;
		16'b0001000010010111 : data_out =  24'b000000000111111101001110;
		16'b0001000010011001 : data_out =  24'b000000000111111101101110;
		16'b0001000010011011 : data_out =  24'b000000000111111110001111;
		16'b0001000010011101 : data_out =  24'b000000000111111110110000;
		16'b0001000010011111 : data_out =  24'b000000000111111111010000;
		16'b0001000010100001 : data_out =  24'b000000000111111111110001;
		16'b0001000010100011 : data_out =  24'b000000001000000000010010;
		16'b0001000010100101 : data_out =  24'b000000001000000000110011;
		16'b0001000010100111 : data_out =  24'b000000001000000001010011;
		16'b0001000010101001 : data_out =  24'b000000001000000001110100;
		16'b0001000010101100 : data_out =  24'b000000001000000010010101;
		16'b0001000010101110 : data_out =  24'b000000001000000010110110;
		16'b0001000010110000 : data_out =  24'b000000001000000011010111;
		16'b0001000010110010 : data_out =  24'b000000001000000011111000;
		16'b0001000010110100 : data_out =  24'b000000001000000100011001;
		16'b0001000010110110 : data_out =  24'b000000001000000100111010;
		16'b0001000010111000 : data_out =  24'b000000001000000101011011;
		16'b0001000010111010 : data_out =  24'b000000001000000101111100;
		16'b0001000010111100 : data_out =  24'b000000001000000110011110;
		16'b0001000010111110 : data_out =  24'b000000001000000110111111;
		16'b0001000011000000 : data_out =  24'b000000001000000111100000;
		16'b0001000011000010 : data_out =  24'b000000001000001000000001;
		16'b0001000011000100 : data_out =  24'b000000001000001000100011;
		16'b0001000011000110 : data_out =  24'b000000001000001001000100;
		16'b0001000011001000 : data_out =  24'b000000001000001001100101;
		16'b0001000011001010 : data_out =  24'b000000001000001010000111;
		16'b0001000011001100 : data_out =  24'b000000001000001010101000;
		16'b0001000011001110 : data_out =  24'b000000001000001011001010;
		16'b0001000011010000 : data_out =  24'b000000001000001011101011;
		16'b0001000011010010 : data_out =  24'b000000001000001100001101;
		16'b0001000011010100 : data_out =  24'b000000001000001100101110;
		16'b0001000011010111 : data_out =  24'b000000001000001101010000;
		16'b0001000011011001 : data_out =  24'b000000001000001101110001;
		16'b0001000011011011 : data_out =  24'b000000001000001110010011;
		16'b0001000011011101 : data_out =  24'b000000001000001110110101;
		16'b0001000011011111 : data_out =  24'b000000001000001111010111;
		16'b0001000011100001 : data_out =  24'b000000001000001111111000;
		16'b0001000011100011 : data_out =  24'b000000001000010000011010;
		16'b0001000011100101 : data_out =  24'b000000001000010000111100;
		16'b0001000011100111 : data_out =  24'b000000001000010001011110;
		16'b0001000011101001 : data_out =  24'b000000001000010010000000;
		16'b0001000011101011 : data_out =  24'b000000001000010010100010;
		16'b0001000011101101 : data_out =  24'b000000001000010011000100;
		16'b0001000011101111 : data_out =  24'b000000001000010011100110;
		16'b0001000011110001 : data_out =  24'b000000001000010100001000;
		16'b0001000011110011 : data_out =  24'b000000001000010100101010;
		16'b0001000011110101 : data_out =  24'b000000001000010101001100;
		16'b0001000011110111 : data_out =  24'b000000001000010101101110;
		16'b0001000011111001 : data_out =  24'b000000001000010110010000;
		16'b0001000011111011 : data_out =  24'b000000001000010110110010;
		16'b0001000011111101 : data_out =  24'b000000001000010111010101;
		16'b0001000011111111 : data_out =  24'b000000001000010111110111;
		16'b0001000100000010 : data_out =  24'b000000001000011000011001;
		16'b0001000100000100 : data_out =  24'b000000001000011000111100;
		16'b0001000100000110 : data_out =  24'b000000001000011001011110;
		16'b0001000100001000 : data_out =  24'b000000001000011010000000;
		16'b0001000100001010 : data_out =  24'b000000001000011010100011;
		16'b0001000100001100 : data_out =  24'b000000001000011011000101;
		16'b0001000100001110 : data_out =  24'b000000001000011011101000;
		16'b0001000100010000 : data_out =  24'b000000001000011100001010;
		16'b0001000100010010 : data_out =  24'b000000001000011100101101;
		16'b0001000100010100 : data_out =  24'b000000001000011101010000;
		16'b0001000100010110 : data_out =  24'b000000001000011101110010;
		16'b0001000100011000 : data_out =  24'b000000001000011110010101;
		16'b0001000100011010 : data_out =  24'b000000001000011110111000;
		16'b0001000100011100 : data_out =  24'b000000001000011111011010;
		16'b0001000100011110 : data_out =  24'b000000001000011111111101;
		16'b0001000100100000 : data_out =  24'b000000001000100000100000;
		16'b0001000100100010 : data_out =  24'b000000001000100001000011;
		16'b0001000100100100 : data_out =  24'b000000001000100001100110;
		16'b0001000100100110 : data_out =  24'b000000001000100010001001;
		16'b0001000100101000 : data_out =  24'b000000001000100010101100;
		16'b0001000100101011 : data_out =  24'b000000001000100011001111;
		16'b0001000100101101 : data_out =  24'b000000001000100011110010;
		16'b0001000100101111 : data_out =  24'b000000001000100100010101;
		16'b0001000100110001 : data_out =  24'b000000001000100100111000;
		16'b0001000100110011 : data_out =  24'b000000001000100101011011;
		16'b0001000100110101 : data_out =  24'b000000001000100101111110;
		16'b0001000100110111 : data_out =  24'b000000001000100110100001;
		16'b0001000100111001 : data_out =  24'b000000001000100111000101;
		16'b0001000100111011 : data_out =  24'b000000001000100111101000;
		16'b0001000100111101 : data_out =  24'b000000001000101000001011;
		16'b0001000100111111 : data_out =  24'b000000001000101000101111;
		16'b0001000101000001 : data_out =  24'b000000001000101001010010;
		16'b0001000101000011 : data_out =  24'b000000001000101001110110;
		16'b0001000101000101 : data_out =  24'b000000001000101010011001;
		16'b0001000101000111 : data_out =  24'b000000001000101010111100;
		16'b0001000101001001 : data_out =  24'b000000001000101011100000;
		16'b0001000101001011 : data_out =  24'b000000001000101100000100;
		16'b0001000101001101 : data_out =  24'b000000001000101100100111;
		16'b0001000101001111 : data_out =  24'b000000001000101101001011;
		16'b0001000101010001 : data_out =  24'b000000001000101101101111;
		16'b0001000101010011 : data_out =  24'b000000001000101110010010;
		16'b0001000101010110 : data_out =  24'b000000001000101110110110;
		16'b0001000101011000 : data_out =  24'b000000001000101111011010;
		16'b0001000101011010 : data_out =  24'b000000001000101111111110;
		16'b0001000101011100 : data_out =  24'b000000001000110000100001;
		16'b0001000101011110 : data_out =  24'b000000001000110001000101;
		16'b0001000101100000 : data_out =  24'b000000001000110001101001;
		16'b0001000101100010 : data_out =  24'b000000001000110010001101;
		16'b0001000101100100 : data_out =  24'b000000001000110010110001;
		16'b0001000101100110 : data_out =  24'b000000001000110011010101;
		16'b0001000101101000 : data_out =  24'b000000001000110011111001;
		16'b0001000101101010 : data_out =  24'b000000001000110100011101;
		16'b0001000101101100 : data_out =  24'b000000001000110101000010;
		16'b0001000101101110 : data_out =  24'b000000001000110101100110;
		16'b0001000101110000 : data_out =  24'b000000001000110110001010;
		16'b0001000101110010 : data_out =  24'b000000001000110110101110;
		16'b0001000101110100 : data_out =  24'b000000001000110111010011;
		16'b0001000101110110 : data_out =  24'b000000001000110111110111;
		16'b0001000101111000 : data_out =  24'b000000001000111000011011;
		16'b0001000101111010 : data_out =  24'b000000001000111001000000;
		16'b0001000101111100 : data_out =  24'b000000001000111001100100;
		16'b0001000101111110 : data_out =  24'b000000001000111010001001;
		16'b0001000110000001 : data_out =  24'b000000001000111010101101;
		16'b0001000110000011 : data_out =  24'b000000001000111011010010;
		16'b0001000110000101 : data_out =  24'b000000001000111011110110;
		16'b0001000110000111 : data_out =  24'b000000001000111100011011;
		16'b0001000110001001 : data_out =  24'b000000001000111100111111;
		16'b0001000110001011 : data_out =  24'b000000001000111101100100;
		16'b0001000110001101 : data_out =  24'b000000001000111110001001;
		16'b0001000110001111 : data_out =  24'b000000001000111110101110;
		16'b0001000110010001 : data_out =  24'b000000001000111111010010;
		16'b0001000110010011 : data_out =  24'b000000001000111111110111;
		16'b0001000110010101 : data_out =  24'b000000001001000000011100;
		16'b0001000110010111 : data_out =  24'b000000001001000001000001;
		16'b0001000110011001 : data_out =  24'b000000001001000001100110;
		16'b0001000110011011 : data_out =  24'b000000001001000010001011;
		16'b0001000110011101 : data_out =  24'b000000001001000010110000;
		16'b0001000110011111 : data_out =  24'b000000001001000011010101;
		16'b0001000110100001 : data_out =  24'b000000001001000011111010;
		16'b0001000110100011 : data_out =  24'b000000001001000100011111;
		16'b0001000110100101 : data_out =  24'b000000001001000101000100;
		16'b0001000110100111 : data_out =  24'b000000001001000101101010;
		16'b0001000110101001 : data_out =  24'b000000001001000110001111;
		16'b0001000110101100 : data_out =  24'b000000001001000110110100;
		16'b0001000110101110 : data_out =  24'b000000001001000111011001;
		16'b0001000110110000 : data_out =  24'b000000001001000111111111;
		16'b0001000110110010 : data_out =  24'b000000001001001000100100;
		16'b0001000110110100 : data_out =  24'b000000001001001001001010;
		16'b0001000110110110 : data_out =  24'b000000001001001001101111;
		16'b0001000110111000 : data_out =  24'b000000001001001010010101;
		16'b0001000110111010 : data_out =  24'b000000001001001010111010;
		16'b0001000110111100 : data_out =  24'b000000001001001011100000;
		16'b0001000110111110 : data_out =  24'b000000001001001100000101;
		16'b0001000111000000 : data_out =  24'b000000001001001100101011;
		16'b0001000111000010 : data_out =  24'b000000001001001101010001;
		16'b0001000111000100 : data_out =  24'b000000001001001101110110;
		16'b0001000111000110 : data_out =  24'b000000001001001110011100;
		16'b0001000111001000 : data_out =  24'b000000001001001111000010;
		16'b0001000111001010 : data_out =  24'b000000001001001111101000;
		16'b0001000111001100 : data_out =  24'b000000001001010000001110;
		16'b0001000111001110 : data_out =  24'b000000001001010000110100;
		16'b0001000111010000 : data_out =  24'b000000001001010001011010;
		16'b0001000111010010 : data_out =  24'b000000001001010010000000;
		16'b0001000111010100 : data_out =  24'b000000001001010010100110;
		16'b0001000111010111 : data_out =  24'b000000001001010011001100;
		16'b0001000111011001 : data_out =  24'b000000001001010011110010;
		16'b0001000111011011 : data_out =  24'b000000001001010100011000;
		16'b0001000111011101 : data_out =  24'b000000001001010100111110;
		16'b0001000111011111 : data_out =  24'b000000001001010101100100;
		16'b0001000111100001 : data_out =  24'b000000001001010110001011;
		16'b0001000111100011 : data_out =  24'b000000001001010110110001;
		16'b0001000111100101 : data_out =  24'b000000001001010111010111;
		16'b0001000111100111 : data_out =  24'b000000001001010111111110;
		16'b0001000111101001 : data_out =  24'b000000001001011000100100;
		16'b0001000111101011 : data_out =  24'b000000001001011001001011;
		16'b0001000111101101 : data_out =  24'b000000001001011001110001;
		16'b0001000111101111 : data_out =  24'b000000001001011010011000;
		16'b0001000111110001 : data_out =  24'b000000001001011010111110;
		16'b0001000111110011 : data_out =  24'b000000001001011011100101;
		16'b0001000111110101 : data_out =  24'b000000001001011100001011;
		16'b0001000111110111 : data_out =  24'b000000001001011100110010;
		16'b0001000111111001 : data_out =  24'b000000001001011101011001;
		16'b0001000111111011 : data_out =  24'b000000001001011110000000;
		16'b0001000111111101 : data_out =  24'b000000001001011110100110;
		16'b0001000111111111 : data_out =  24'b000000001001011111001101;
		16'b0001001000000010 : data_out =  24'b000000001001011111110100;
		16'b0001001000000100 : data_out =  24'b000000001001100000011011;
		16'b0001001000000110 : data_out =  24'b000000001001100001000010;
		16'b0001001000001000 : data_out =  24'b000000001001100001101001;
		16'b0001001000001010 : data_out =  24'b000000001001100010010000;
		16'b0001001000001100 : data_out =  24'b000000001001100010110111;
		16'b0001001000001110 : data_out =  24'b000000001001100011011110;
		16'b0001001000010000 : data_out =  24'b000000001001100100000101;
		16'b0001001000010010 : data_out =  24'b000000001001100100101101;
		16'b0001001000010100 : data_out =  24'b000000001001100101010100;
		16'b0001001000010110 : data_out =  24'b000000001001100101111011;
		16'b0001001000011000 : data_out =  24'b000000001001100110100010;
		16'b0001001000011010 : data_out =  24'b000000001001100111001010;
		16'b0001001000011100 : data_out =  24'b000000001001100111110001;
		16'b0001001000011110 : data_out =  24'b000000001001101000011001;
		16'b0001001000100000 : data_out =  24'b000000001001101001000000;
		16'b0001001000100010 : data_out =  24'b000000001001101001101000;
		16'b0001001000100100 : data_out =  24'b000000001001101010001111;
		16'b0001001000100110 : data_out =  24'b000000001001101010110111;
		16'b0001001000101000 : data_out =  24'b000000001001101011011110;
		16'b0001001000101011 : data_out =  24'b000000001001101100000110;
		16'b0001001000101101 : data_out =  24'b000000001001101100101110;
		16'b0001001000101111 : data_out =  24'b000000001001101101010101;
		16'b0001001000110001 : data_out =  24'b000000001001101101111101;
		16'b0001001000110011 : data_out =  24'b000000001001101110100101;
		16'b0001001000110101 : data_out =  24'b000000001001101111001101;
		16'b0001001000110111 : data_out =  24'b000000001001101111110101;
		16'b0001001000111001 : data_out =  24'b000000001001110000011101;
		16'b0001001000111011 : data_out =  24'b000000001001110001000101;
		16'b0001001000111101 : data_out =  24'b000000001001110001101101;
		16'b0001001000111111 : data_out =  24'b000000001001110010010101;
		16'b0001001001000001 : data_out =  24'b000000001001110010111101;
		16'b0001001001000011 : data_out =  24'b000000001001110011100101;
		16'b0001001001000101 : data_out =  24'b000000001001110100001101;
		16'b0001001001000111 : data_out =  24'b000000001001110100110110;
		16'b0001001001001001 : data_out =  24'b000000001001110101011110;
		16'b0001001001001011 : data_out =  24'b000000001001110110000110;
		16'b0001001001001101 : data_out =  24'b000000001001110110101110;
		16'b0001001001001111 : data_out =  24'b000000001001110111010111;
		16'b0001001001010001 : data_out =  24'b000000001001110111111111;
		16'b0001001001010011 : data_out =  24'b000000001001111000101000;
		16'b0001001001010110 : data_out =  24'b000000001001111001010000;
		16'b0001001001011000 : data_out =  24'b000000001001111001111001;
		16'b0001001001011010 : data_out =  24'b000000001001111010100001;
		16'b0001001001011100 : data_out =  24'b000000001001111011001010;
		16'b0001001001011110 : data_out =  24'b000000001001111011110011;
		16'b0001001001100000 : data_out =  24'b000000001001111100011011;
		16'b0001001001100010 : data_out =  24'b000000001001111101000100;
		16'b0001001001100100 : data_out =  24'b000000001001111101101101;
		16'b0001001001100110 : data_out =  24'b000000001001111110010110;
		16'b0001001001101000 : data_out =  24'b000000001001111110111111;
		16'b0001001001101010 : data_out =  24'b000000001001111111101000;
		16'b0001001001101100 : data_out =  24'b000000001010000000010000;
		16'b0001001001101110 : data_out =  24'b000000001010000000111001;
		16'b0001001001110000 : data_out =  24'b000000001010000001100011;
		16'b0001001001110010 : data_out =  24'b000000001010000010001100;
		16'b0001001001110100 : data_out =  24'b000000001010000010110101;
		16'b0001001001110110 : data_out =  24'b000000001010000011011110;
		16'b0001001001111000 : data_out =  24'b000000001010000100000111;
		16'b0001001001111010 : data_out =  24'b000000001010000100110000;
		16'b0001001001111100 : data_out =  24'b000000001010000101011010;
		16'b0001001001111110 : data_out =  24'b000000001010000110000011;
		16'b0001001010000001 : data_out =  24'b000000001010000110101100;
		16'b0001001010000011 : data_out =  24'b000000001010000111010110;
		16'b0001001010000101 : data_out =  24'b000000001010000111111111;
		16'b0001001010000111 : data_out =  24'b000000001010001000101001;
		16'b0001001010001001 : data_out =  24'b000000001010001001010010;
		16'b0001001010001011 : data_out =  24'b000000001010001001111100;
		16'b0001001010001101 : data_out =  24'b000000001010001010100101;
		16'b0001001010001111 : data_out =  24'b000000001010001011001111;
		16'b0001001010010001 : data_out =  24'b000000001010001011111001;
		16'b0001001010010011 : data_out =  24'b000000001010001100100011;
		16'b0001001010010101 : data_out =  24'b000000001010001101001100;
		16'b0001001010010111 : data_out =  24'b000000001010001101110110;
		16'b0001001010011001 : data_out =  24'b000000001010001110100000;
		16'b0001001010011011 : data_out =  24'b000000001010001111001010;
		16'b0001001010011101 : data_out =  24'b000000001010001111110100;
		16'b0001001010011111 : data_out =  24'b000000001010010000011110;
		16'b0001001010100001 : data_out =  24'b000000001010010001001000;
		16'b0001001010100011 : data_out =  24'b000000001010010001110010;
		16'b0001001010100101 : data_out =  24'b000000001010010010011100;
		16'b0001001010100111 : data_out =  24'b000000001010010011000110;
		16'b0001001010101001 : data_out =  24'b000000001010010011110000;
		16'b0001001010101100 : data_out =  24'b000000001010010100011011;
		16'b0001001010101110 : data_out =  24'b000000001010010101000101;
		16'b0001001010110000 : data_out =  24'b000000001010010101101111;
		16'b0001001010110010 : data_out =  24'b000000001010010110011010;
		16'b0001001010110100 : data_out =  24'b000000001010010111000100;
		16'b0001001010110110 : data_out =  24'b000000001010010111101111;
		16'b0001001010111000 : data_out =  24'b000000001010011000011001;
		16'b0001001010111010 : data_out =  24'b000000001010011001000100;
		16'b0001001010111100 : data_out =  24'b000000001010011001101110;
		16'b0001001010111110 : data_out =  24'b000000001010011010011001;
		16'b0001001011000000 : data_out =  24'b000000001010011011000011;
		16'b0001001011000010 : data_out =  24'b000000001010011011101110;
		16'b0001001011000100 : data_out =  24'b000000001010011100011001;
		16'b0001001011000110 : data_out =  24'b000000001010011101000100;
		16'b0001001011001000 : data_out =  24'b000000001010011101101111;
		16'b0001001011001010 : data_out =  24'b000000001010011110011001;
		16'b0001001011001100 : data_out =  24'b000000001010011111000100;
		16'b0001001011001110 : data_out =  24'b000000001010011111101111;
		16'b0001001011010000 : data_out =  24'b000000001010100000011010;
		16'b0001001011010010 : data_out =  24'b000000001010100001000101;
		16'b0001001011010100 : data_out =  24'b000000001010100001110001;
		16'b0001001011010111 : data_out =  24'b000000001010100010011100;
		16'b0001001011011001 : data_out =  24'b000000001010100011000111;
		16'b0001001011011011 : data_out =  24'b000000001010100011110010;
		16'b0001001011011101 : data_out =  24'b000000001010100100011101;
		16'b0001001011011111 : data_out =  24'b000000001010100101001001;
		16'b0001001011100001 : data_out =  24'b000000001010100101110100;
		16'b0001001011100011 : data_out =  24'b000000001010100110011111;
		16'b0001001011100101 : data_out =  24'b000000001010100111001011;
		16'b0001001011100111 : data_out =  24'b000000001010100111110110;
		16'b0001001011101001 : data_out =  24'b000000001010101000100010;
		16'b0001001011101011 : data_out =  24'b000000001010101001001101;
		16'b0001001011101101 : data_out =  24'b000000001010101001111001;
		16'b0001001011101111 : data_out =  24'b000000001010101010100101;
		16'b0001001011110001 : data_out =  24'b000000001010101011010000;
		16'b0001001011110011 : data_out =  24'b000000001010101011111100;
		16'b0001001011110101 : data_out =  24'b000000001010101100101000;
		16'b0001001011110111 : data_out =  24'b000000001010101101010100;
		16'b0001001011111001 : data_out =  24'b000000001010101110000000;
		16'b0001001011111011 : data_out =  24'b000000001010101110101100;
		16'b0001001011111101 : data_out =  24'b000000001010101111011000;
		16'b0001001011111111 : data_out =  24'b000000001010110000000100;
		16'b0001001100000010 : data_out =  24'b000000001010110000110000;
		16'b0001001100000100 : data_out =  24'b000000001010110001011100;
		16'b0001001100000110 : data_out =  24'b000000001010110010001000;
		16'b0001001100001000 : data_out =  24'b000000001010110010110100;
		16'b0001001100001010 : data_out =  24'b000000001010110011100000;
		16'b0001001100001100 : data_out =  24'b000000001010110100001101;
		16'b0001001100001110 : data_out =  24'b000000001010110100111001;
		16'b0001001100010000 : data_out =  24'b000000001010110101100101;
		16'b0001001100010010 : data_out =  24'b000000001010110110010010;
		16'b0001001100010100 : data_out =  24'b000000001010110110111110;
		16'b0001001100010110 : data_out =  24'b000000001010110111101011;
		16'b0001001100011000 : data_out =  24'b000000001010111000010111;
		16'b0001001100011010 : data_out =  24'b000000001010111001000100;
		16'b0001001100011100 : data_out =  24'b000000001010111001110000;
		16'b0001001100011110 : data_out =  24'b000000001010111010011101;
		16'b0001001100100000 : data_out =  24'b000000001010111011001010;
		16'b0001001100100010 : data_out =  24'b000000001010111011110111;
		16'b0001001100100100 : data_out =  24'b000000001010111100100011;
		16'b0001001100100110 : data_out =  24'b000000001010111101010000;
		16'b0001001100101000 : data_out =  24'b000000001010111101111101;
		16'b0001001100101011 : data_out =  24'b000000001010111110101010;
		16'b0001001100101101 : data_out =  24'b000000001010111111010111;
		16'b0001001100101111 : data_out =  24'b000000001011000000000100;
		16'b0001001100110001 : data_out =  24'b000000001011000000110001;
		16'b0001001100110011 : data_out =  24'b000000001011000001011110;
		16'b0001001100110101 : data_out =  24'b000000001011000010001100;
		16'b0001001100110111 : data_out =  24'b000000001011000010111001;
		16'b0001001100111001 : data_out =  24'b000000001011000011100110;
		16'b0001001100111011 : data_out =  24'b000000001011000100010011;
		16'b0001001100111101 : data_out =  24'b000000001011000101000001;
		16'b0001001100111111 : data_out =  24'b000000001011000101101110;
		16'b0001001101000001 : data_out =  24'b000000001011000110011100;
		16'b0001001101000011 : data_out =  24'b000000001011000111001001;
		16'b0001001101000101 : data_out =  24'b000000001011000111110111;
		16'b0001001101000111 : data_out =  24'b000000001011001000100100;
		16'b0001001101001001 : data_out =  24'b000000001011001001010010;
		16'b0001001101001011 : data_out =  24'b000000001011001010000000;
		16'b0001001101001101 : data_out =  24'b000000001011001010101101;
		16'b0001001101001111 : data_out =  24'b000000001011001011011011;
		16'b0001001101010001 : data_out =  24'b000000001011001100001001;
		16'b0001001101010011 : data_out =  24'b000000001011001100110111;
		16'b0001001101010110 : data_out =  24'b000000001011001101100101;
		16'b0001001101011000 : data_out =  24'b000000001011001110010011;
		16'b0001001101011010 : data_out =  24'b000000001011001111000000;
		16'b0001001101011100 : data_out =  24'b000000001011001111101111;
		16'b0001001101011110 : data_out =  24'b000000001011010000011101;
		16'b0001001101100000 : data_out =  24'b000000001011010001001011;
		16'b0001001101100010 : data_out =  24'b000000001011010001111001;
		16'b0001001101100100 : data_out =  24'b000000001011010010100111;
		16'b0001001101100110 : data_out =  24'b000000001011010011010101;
		16'b0001001101101000 : data_out =  24'b000000001011010100000100;
		16'b0001001101101010 : data_out =  24'b000000001011010100110010;
		16'b0001001101101100 : data_out =  24'b000000001011010101100001;
		16'b0001001101101110 : data_out =  24'b000000001011010110001111;
		16'b0001001101110000 : data_out =  24'b000000001011010110111101;
		16'b0001001101110010 : data_out =  24'b000000001011010111101100;
		16'b0001001101110100 : data_out =  24'b000000001011011000011011;
		16'b0001001101110110 : data_out =  24'b000000001011011001001001;
		16'b0001001101111000 : data_out =  24'b000000001011011001111000;
		16'b0001001101111010 : data_out =  24'b000000001011011010100111;
		16'b0001001101111100 : data_out =  24'b000000001011011011010101;
		16'b0001001101111110 : data_out =  24'b000000001011011100000100;
		16'b0001001110000001 : data_out =  24'b000000001011011100110011;
		16'b0001001110000011 : data_out =  24'b000000001011011101100010;
		16'b0001001110000101 : data_out =  24'b000000001011011110010001;
		16'b0001001110000111 : data_out =  24'b000000001011011111000000;
		16'b0001001110001001 : data_out =  24'b000000001011011111101111;
		16'b0001001110001011 : data_out =  24'b000000001011100000011110;
		16'b0001001110001101 : data_out =  24'b000000001011100001001101;
		16'b0001001110001111 : data_out =  24'b000000001011100001111101;
		16'b0001001110010001 : data_out =  24'b000000001011100010101100;
		16'b0001001110010011 : data_out =  24'b000000001011100011011011;
		16'b0001001110010101 : data_out =  24'b000000001011100100001011;
		16'b0001001110010111 : data_out =  24'b000000001011100100111010;
		16'b0001001110011001 : data_out =  24'b000000001011100101101001;
		16'b0001001110011011 : data_out =  24'b000000001011100110011001;
		16'b0001001110011101 : data_out =  24'b000000001011100111001000;
		16'b0001001110011111 : data_out =  24'b000000001011100111111000;
		16'b0001001110100001 : data_out =  24'b000000001011101000101000;
		16'b0001001110100011 : data_out =  24'b000000001011101001010111;
		16'b0001001110100101 : data_out =  24'b000000001011101010000111;
		16'b0001001110100111 : data_out =  24'b000000001011101010110111;
		16'b0001001110101001 : data_out =  24'b000000001011101011100111;
		16'b0001001110101100 : data_out =  24'b000000001011101100010110;
		16'b0001001110101110 : data_out =  24'b000000001011101101000110;
		16'b0001001110110000 : data_out =  24'b000000001011101101110110;
		16'b0001001110110010 : data_out =  24'b000000001011101110100110;
		16'b0001001110110100 : data_out =  24'b000000001011101111010110;
		16'b0001001110110110 : data_out =  24'b000000001011110000000111;
		16'b0001001110111000 : data_out =  24'b000000001011110000110111;
		16'b0001001110111010 : data_out =  24'b000000001011110001100111;
		16'b0001001110111100 : data_out =  24'b000000001011110010010111;
		16'b0001001110111110 : data_out =  24'b000000001011110011000111;
		16'b0001001111000000 : data_out =  24'b000000001011110011111000;
		16'b0001001111000010 : data_out =  24'b000000001011110100101000;
		16'b0001001111000100 : data_out =  24'b000000001011110101011001;
		16'b0001001111000110 : data_out =  24'b000000001011110110001001;
		16'b0001001111001000 : data_out =  24'b000000001011110110111010;
		16'b0001001111001010 : data_out =  24'b000000001011110111101010;
		16'b0001001111001100 : data_out =  24'b000000001011111000011011;
		16'b0001001111001110 : data_out =  24'b000000001011111001001100;
		16'b0001001111010000 : data_out =  24'b000000001011111001111100;
		16'b0001001111010010 : data_out =  24'b000000001011111010101101;
		16'b0001001111010100 : data_out =  24'b000000001011111011011110;
		16'b0001001111010111 : data_out =  24'b000000001011111100001111;
		16'b0001001111011001 : data_out =  24'b000000001011111101000000;
		16'b0001001111011011 : data_out =  24'b000000001011111101110001;
		16'b0001001111011101 : data_out =  24'b000000001011111110100010;
		16'b0001001111011111 : data_out =  24'b000000001011111111010011;
		16'b0001001111100001 : data_out =  24'b000000001100000000000100;
		16'b0001001111100011 : data_out =  24'b000000001100000000110101;
		16'b0001001111100101 : data_out =  24'b000000001100000001100111;
		16'b0001001111100111 : data_out =  24'b000000001100000010011000;
		16'b0001001111101001 : data_out =  24'b000000001100000011001001;
		16'b0001001111101011 : data_out =  24'b000000001100000011111010;
		16'b0001001111101101 : data_out =  24'b000000001100000100101100;
		16'b0001001111101111 : data_out =  24'b000000001100000101011101;
		16'b0001001111110001 : data_out =  24'b000000001100000110001111;
		16'b0001001111110011 : data_out =  24'b000000001100000111000000;
		16'b0001001111110101 : data_out =  24'b000000001100000111110010;
		16'b0001001111110111 : data_out =  24'b000000001100001000100100;
		16'b0001001111111001 : data_out =  24'b000000001100001001010110;
		16'b0001001111111011 : data_out =  24'b000000001100001010000111;
		16'b0001001111111101 : data_out =  24'b000000001100001010111001;
		16'b0001001111111111 : data_out =  24'b000000001100001011101011;
		16'b0001010000000010 : data_out =  24'b000000001100001100011101;
		16'b0001010000000100 : data_out =  24'b000000001100001101001111;
		16'b0001010000000110 : data_out =  24'b000000001100001110000001;
		16'b0001010000001000 : data_out =  24'b000000001100001110110011;
		16'b0001010000001010 : data_out =  24'b000000001100001111100101;
		16'b0001010000001100 : data_out =  24'b000000001100010000010111;
		16'b0001010000001110 : data_out =  24'b000000001100010001001010;
		16'b0001010000010000 : data_out =  24'b000000001100010001111100;
		16'b0001010000010010 : data_out =  24'b000000001100010010101110;
		16'b0001010000010100 : data_out =  24'b000000001100010011100000;
		16'b0001010000010110 : data_out =  24'b000000001100010100010011;
		16'b0001010000011000 : data_out =  24'b000000001100010101000101;
		16'b0001010000011010 : data_out =  24'b000000001100010101111000;
		16'b0001010000011100 : data_out =  24'b000000001100010110101011;
		16'b0001010000011110 : data_out =  24'b000000001100010111011101;
		16'b0001010000100000 : data_out =  24'b000000001100011000010000;
		16'b0001010000100010 : data_out =  24'b000000001100011001000011;
		16'b0001010000100100 : data_out =  24'b000000001100011001110101;
		16'b0001010000100110 : data_out =  24'b000000001100011010101000;
		16'b0001010000101000 : data_out =  24'b000000001100011011011011;
		16'b0001010000101011 : data_out =  24'b000000001100011100001110;
		16'b0001010000101101 : data_out =  24'b000000001100011101000001;
		16'b0001010000101111 : data_out =  24'b000000001100011101110100;
		16'b0001010000110001 : data_out =  24'b000000001100011110100111;
		16'b0001010000110011 : data_out =  24'b000000001100011111011010;
		16'b0001010000110101 : data_out =  24'b000000001100100000001101;
		16'b0001010000110111 : data_out =  24'b000000001100100001000001;
		16'b0001010000111001 : data_out =  24'b000000001100100001110100;
		16'b0001010000111011 : data_out =  24'b000000001100100010100111;
		16'b0001010000111101 : data_out =  24'b000000001100100011011011;
		16'b0001010000111111 : data_out =  24'b000000001100100100001110;
		16'b0001010001000001 : data_out =  24'b000000001100100101000010;
		16'b0001010001000011 : data_out =  24'b000000001100100101110101;
		16'b0001010001000101 : data_out =  24'b000000001100100110101001;
		16'b0001010001000111 : data_out =  24'b000000001100100111011100;
		16'b0001010001001001 : data_out =  24'b000000001100101000010000;
		16'b0001010001001011 : data_out =  24'b000000001100101001000100;
		16'b0001010001001101 : data_out =  24'b000000001100101001111000;
		16'b0001010001001111 : data_out =  24'b000000001100101010101100;
		16'b0001010001010001 : data_out =  24'b000000001100101011011111;
		16'b0001010001010011 : data_out =  24'b000000001100101100010011;
		16'b0001010001010110 : data_out =  24'b000000001100101101000111;
		16'b0001010001011000 : data_out =  24'b000000001100101101111011;
		16'b0001010001011010 : data_out =  24'b000000001100101110110000;
		16'b0001010001011100 : data_out =  24'b000000001100101111100100;
		16'b0001010001011110 : data_out =  24'b000000001100110000011000;
		16'b0001010001100000 : data_out =  24'b000000001100110001001100;
		16'b0001010001100010 : data_out =  24'b000000001100110010000001;
		16'b0001010001100100 : data_out =  24'b000000001100110010110101;
		16'b0001010001100110 : data_out =  24'b000000001100110011101001;
		16'b0001010001101000 : data_out =  24'b000000001100110100011110;
		16'b0001010001101010 : data_out =  24'b000000001100110101010010;
		16'b0001010001101100 : data_out =  24'b000000001100110110000111;
		16'b0001010001101110 : data_out =  24'b000000001100110110111100;
		16'b0001010001110000 : data_out =  24'b000000001100110111110000;
		16'b0001010001110010 : data_out =  24'b000000001100111000100101;
		16'b0001010001110100 : data_out =  24'b000000001100111001011010;
		16'b0001010001110110 : data_out =  24'b000000001100111010001111;
		16'b0001010001111000 : data_out =  24'b000000001100111011000100;
		16'b0001010001111010 : data_out =  24'b000000001100111011111001;
		16'b0001010001111100 : data_out =  24'b000000001100111100101110;
		16'b0001010001111110 : data_out =  24'b000000001100111101100011;
		16'b0001010010000001 : data_out =  24'b000000001100111110011000;
		16'b0001010010000011 : data_out =  24'b000000001100111111001101;
		16'b0001010010000101 : data_out =  24'b000000001101000000000010;
		16'b0001010010000111 : data_out =  24'b000000001101000000110111;
		16'b0001010010001001 : data_out =  24'b000000001101000001101101;
		16'b0001010010001011 : data_out =  24'b000000001101000010100010;
		16'b0001010010001101 : data_out =  24'b000000001101000011011000;
		16'b0001010010001111 : data_out =  24'b000000001101000100001101;
		16'b0001010010010001 : data_out =  24'b000000001101000101000011;
		16'b0001010010010011 : data_out =  24'b000000001101000101111000;
		16'b0001010010010101 : data_out =  24'b000000001101000110101110;
		16'b0001010010010111 : data_out =  24'b000000001101000111100100;
		16'b0001010010011001 : data_out =  24'b000000001101001000011001;
		16'b0001010010011011 : data_out =  24'b000000001101001001001111;
		16'b0001010010011101 : data_out =  24'b000000001101001010000101;
		16'b0001010010011111 : data_out =  24'b000000001101001010111011;
		16'b0001010010100001 : data_out =  24'b000000001101001011110001;
		16'b0001010010100011 : data_out =  24'b000000001101001100100111;
		16'b0001010010100101 : data_out =  24'b000000001101001101011101;
		16'b0001010010100111 : data_out =  24'b000000001101001110010011;
		16'b0001010010101001 : data_out =  24'b000000001101001111001001;
		16'b0001010010101100 : data_out =  24'b000000001101010000000000;
		16'b0001010010101110 : data_out =  24'b000000001101010000110110;
		16'b0001010010110000 : data_out =  24'b000000001101010001101100;
		16'b0001010010110010 : data_out =  24'b000000001101010010100011;
		16'b0001010010110100 : data_out =  24'b000000001101010011011001;
		16'b0001010010110110 : data_out =  24'b000000001101010100010000;
		16'b0001010010111000 : data_out =  24'b000000001101010101000110;
		16'b0001010010111010 : data_out =  24'b000000001101010101111101;
		16'b0001010010111100 : data_out =  24'b000000001101010110110100;
		16'b0001010010111110 : data_out =  24'b000000001101010111101010;
		16'b0001010011000000 : data_out =  24'b000000001101011000100001;
		16'b0001010011000010 : data_out =  24'b000000001101011001011000;
		16'b0001010011000100 : data_out =  24'b000000001101011010001111;
		16'b0001010011000110 : data_out =  24'b000000001101011011000110;
		16'b0001010011001000 : data_out =  24'b000000001101011011111101;
		16'b0001010011001010 : data_out =  24'b000000001101011100110100;
		16'b0001010011001100 : data_out =  24'b000000001101011101101011;
		16'b0001010011001110 : data_out =  24'b000000001101011110100010;
		16'b0001010011010000 : data_out =  24'b000000001101011111011001;
		16'b0001010011010010 : data_out =  24'b000000001101100000010001;
		16'b0001010011010100 : data_out =  24'b000000001101100001001000;
		16'b0001010011010111 : data_out =  24'b000000001101100001111111;
		16'b0001010011011001 : data_out =  24'b000000001101100010110111;
		16'b0001010011011011 : data_out =  24'b000000001101100011101110;
		16'b0001010011011101 : data_out =  24'b000000001101100100100110;
		16'b0001010011011111 : data_out =  24'b000000001101100101011110;
		16'b0001010011100001 : data_out =  24'b000000001101100110010101;
		16'b0001010011100011 : data_out =  24'b000000001101100111001101;
		16'b0001010011100101 : data_out =  24'b000000001101101000000101;
		16'b0001010011100111 : data_out =  24'b000000001101101000111101;
		16'b0001010011101001 : data_out =  24'b000000001101101001110100;
		16'b0001010011101011 : data_out =  24'b000000001101101010101100;
		16'b0001010011101101 : data_out =  24'b000000001101101011100100;
		16'b0001010011101111 : data_out =  24'b000000001101101100011100;
		16'b0001010011110001 : data_out =  24'b000000001101101101010101;
		16'b0001010011110011 : data_out =  24'b000000001101101110001101;
		16'b0001010011110101 : data_out =  24'b000000001101101111000101;
		16'b0001010011110111 : data_out =  24'b000000001101101111111101;
		16'b0001010011111001 : data_out =  24'b000000001101110000110110;
		16'b0001010011111011 : data_out =  24'b000000001101110001101110;
		16'b0001010011111101 : data_out =  24'b000000001101110010100111;
		16'b0001010011111111 : data_out =  24'b000000001101110011011111;
		16'b0001010100000010 : data_out =  24'b000000001101110100011000;
		16'b0001010100000100 : data_out =  24'b000000001101110101010000;
		16'b0001010100000110 : data_out =  24'b000000001101110110001001;
		16'b0001010100001000 : data_out =  24'b000000001101110111000010;
		16'b0001010100001010 : data_out =  24'b000000001101110111111010;
		16'b0001010100001100 : data_out =  24'b000000001101111000110011;
		16'b0001010100001110 : data_out =  24'b000000001101111001101100;
		16'b0001010100010000 : data_out =  24'b000000001101111010100101;
		16'b0001010100010010 : data_out =  24'b000000001101111011011110;
		16'b0001010100010100 : data_out =  24'b000000001101111100010111;
		16'b0001010100010110 : data_out =  24'b000000001101111101010000;
		16'b0001010100011000 : data_out =  24'b000000001101111110001010;
		16'b0001010100011010 : data_out =  24'b000000001101111111000011;
		16'b0001010100011100 : data_out =  24'b000000001101111111111100;
		16'b0001010100011110 : data_out =  24'b000000001110000000110110;
		16'b0001010100100000 : data_out =  24'b000000001110000001101111;
		16'b0001010100100010 : data_out =  24'b000000001110000010101000;
		16'b0001010100100100 : data_out =  24'b000000001110000011100010;
		16'b0001010100100110 : data_out =  24'b000000001110000100011100;
		16'b0001010100101000 : data_out =  24'b000000001110000101010101;
		16'b0001010100101011 : data_out =  24'b000000001110000110001111;
		16'b0001010100101101 : data_out =  24'b000000001110000111001001;
		16'b0001010100101111 : data_out =  24'b000000001110001000000011;
		16'b0001010100110001 : data_out =  24'b000000001110001000111100;
		16'b0001010100110011 : data_out =  24'b000000001110001001110110;
		16'b0001010100110101 : data_out =  24'b000000001110001010110000;
		16'b0001010100110111 : data_out =  24'b000000001110001011101011;
		16'b0001010100111001 : data_out =  24'b000000001110001100100101;
		16'b0001010100111011 : data_out =  24'b000000001110001101011111;
		16'b0001010100111101 : data_out =  24'b000000001110001110011001;
		16'b0001010100111111 : data_out =  24'b000000001110001111010011;
		16'b0001010101000001 : data_out =  24'b000000001110010000001110;
		16'b0001010101000011 : data_out =  24'b000000001110010001001000;
		16'b0001010101000101 : data_out =  24'b000000001110010010000011;
		16'b0001010101000111 : data_out =  24'b000000001110010010111101;
		16'b0001010101001001 : data_out =  24'b000000001110010011111000;
		16'b0001010101001011 : data_out =  24'b000000001110010100110010;
		16'b0001010101001101 : data_out =  24'b000000001110010101101101;
		16'b0001010101001111 : data_out =  24'b000000001110010110101000;
		16'b0001010101010001 : data_out =  24'b000000001110010111100011;
		16'b0001010101010011 : data_out =  24'b000000001110011000011110;
		16'b0001010101010110 : data_out =  24'b000000001110011001011000;
		16'b0001010101011000 : data_out =  24'b000000001110011010010011;
		16'b0001010101011010 : data_out =  24'b000000001110011011001110;
		16'b0001010101011100 : data_out =  24'b000000001110011100001010;
		16'b0001010101011110 : data_out =  24'b000000001110011101000101;
		16'b0001010101100000 : data_out =  24'b000000001110011110000000;
		16'b0001010101100010 : data_out =  24'b000000001110011110111011;
		16'b0001010101100100 : data_out =  24'b000000001110011111110111;
		16'b0001010101100110 : data_out =  24'b000000001110100000110010;
		16'b0001010101101000 : data_out =  24'b000000001110100001101110;
		16'b0001010101101010 : data_out =  24'b000000001110100010101001;
		16'b0001010101101100 : data_out =  24'b000000001110100011100101;
		16'b0001010101101110 : data_out =  24'b000000001110100100100000;
		16'b0001010101110000 : data_out =  24'b000000001110100101011100;
		16'b0001010101110010 : data_out =  24'b000000001110100110011000;
		16'b0001010101110100 : data_out =  24'b000000001110100111010100;
		16'b0001010101110110 : data_out =  24'b000000001110101000010000;
		16'b0001010101111000 : data_out =  24'b000000001110101001001011;
		16'b0001010101111010 : data_out =  24'b000000001110101010000111;
		16'b0001010101111100 : data_out =  24'b000000001110101011000100;
		16'b0001010101111110 : data_out =  24'b000000001110101100000000;
		16'b0001010110000001 : data_out =  24'b000000001110101100111100;
		16'b0001010110000011 : data_out =  24'b000000001110101101111000;
		16'b0001010110000101 : data_out =  24'b000000001110101110110100;
		16'b0001010110000111 : data_out =  24'b000000001110101111110001;
		16'b0001010110001001 : data_out =  24'b000000001110110000101101;
		16'b0001010110001011 : data_out =  24'b000000001110110001101010;
		16'b0001010110001101 : data_out =  24'b000000001110110010100110;
		16'b0001010110001111 : data_out =  24'b000000001110110011100011;
		16'b0001010110010001 : data_out =  24'b000000001110110100100000;
		16'b0001010110010011 : data_out =  24'b000000001110110101011100;
		16'b0001010110010101 : data_out =  24'b000000001110110110011001;
		16'b0001010110010111 : data_out =  24'b000000001110110111010110;
		16'b0001010110011001 : data_out =  24'b000000001110111000010011;
		16'b0001010110011011 : data_out =  24'b000000001110111001010000;
		16'b0001010110011101 : data_out =  24'b000000001110111010001101;
		16'b0001010110011111 : data_out =  24'b000000001110111011001010;
		16'b0001010110100001 : data_out =  24'b000000001110111100000111;
		16'b0001010110100011 : data_out =  24'b000000001110111101000100;
		16'b0001010110100101 : data_out =  24'b000000001110111110000010;
		16'b0001010110100111 : data_out =  24'b000000001110111110111111;
		16'b0001010110101001 : data_out =  24'b000000001110111111111100;
		16'b0001010110101100 : data_out =  24'b000000001111000000111010;
		16'b0001010110101110 : data_out =  24'b000000001111000001110111;
		16'b0001010110110000 : data_out =  24'b000000001111000010110101;
		16'b0001010110110010 : data_out =  24'b000000001111000011110011;
		16'b0001010110110100 : data_out =  24'b000000001111000100110000;
		16'b0001010110110110 : data_out =  24'b000000001111000101101110;
		16'b0001010110111000 : data_out =  24'b000000001111000110101100;
		16'b0001010110111010 : data_out =  24'b000000001111000111101010;
		16'b0001010110111100 : data_out =  24'b000000001111001000101000;
		16'b0001010110111110 : data_out =  24'b000000001111001001100110;
		16'b0001010111000000 : data_out =  24'b000000001111001010100100;
		16'b0001010111000010 : data_out =  24'b000000001111001011100010;
		16'b0001010111000100 : data_out =  24'b000000001111001100100000;
		16'b0001010111000110 : data_out =  24'b000000001111001101011111;
		16'b0001010111001000 : data_out =  24'b000000001111001110011101;
		16'b0001010111001010 : data_out =  24'b000000001111001111011011;
		16'b0001010111001100 : data_out =  24'b000000001111010000011010;
		16'b0001010111001110 : data_out =  24'b000000001111010001011000;
		16'b0001010111010000 : data_out =  24'b000000001111010010010111;
		16'b0001010111010010 : data_out =  24'b000000001111010011010110;
		16'b0001010111010100 : data_out =  24'b000000001111010100010100;
		16'b0001010111010111 : data_out =  24'b000000001111010101010011;
		16'b0001010111011001 : data_out =  24'b000000001111010110010010;
		16'b0001010111011011 : data_out =  24'b000000001111010111010001;
		16'b0001010111011101 : data_out =  24'b000000001111011000010000;
		16'b0001010111011111 : data_out =  24'b000000001111011001001111;
		16'b0001010111100001 : data_out =  24'b000000001111011010001110;
		16'b0001010111100011 : data_out =  24'b000000001111011011001101;
		16'b0001010111100101 : data_out =  24'b000000001111011100001100;
		16'b0001010111100111 : data_out =  24'b000000001111011101001011;
		16'b0001010111101001 : data_out =  24'b000000001111011110001011;
		16'b0001010111101011 : data_out =  24'b000000001111011111001010;
		16'b0001010111101101 : data_out =  24'b000000001111100000001010;
		16'b0001010111101111 : data_out =  24'b000000001111100001001001;
		16'b0001010111110001 : data_out =  24'b000000001111100010001001;
		16'b0001010111110011 : data_out =  24'b000000001111100011001000;
		16'b0001010111110101 : data_out =  24'b000000001111100100001000;
		16'b0001010111110111 : data_out =  24'b000000001111100101001000;
		16'b0001010111111001 : data_out =  24'b000000001111100110001000;
		16'b0001010111111011 : data_out =  24'b000000001111100111001000;
		16'b0001010111111101 : data_out =  24'b000000001111101000001000;
		16'b0001010111111111 : data_out =  24'b000000001111101001001000;
		16'b0001011000000010 : data_out =  24'b000000001111101010001000;
		16'b0001011000000100 : data_out =  24'b000000001111101011001000;
		16'b0001011000000110 : data_out =  24'b000000001111101100001000;
		16'b0001011000001000 : data_out =  24'b000000001111101101001001;
		16'b0001011000001010 : data_out =  24'b000000001111101110001001;
		16'b0001011000001100 : data_out =  24'b000000001111101111001001;
		16'b0001011000001110 : data_out =  24'b000000001111110000001010;
		16'b0001011000010000 : data_out =  24'b000000001111110001001010;
		16'b0001011000010010 : data_out =  24'b000000001111110010001011;
		16'b0001011000010100 : data_out =  24'b000000001111110011001100;
		16'b0001011000010110 : data_out =  24'b000000001111110100001100;
		16'b0001011000011000 : data_out =  24'b000000001111110101001101;
		16'b0001011000011010 : data_out =  24'b000000001111110110001110;
		16'b0001011000011100 : data_out =  24'b000000001111110111001111;
		16'b0001011000011110 : data_out =  24'b000000001111111000010000;
		16'b0001011000100000 : data_out =  24'b000000001111111001010001;
		16'b0001011000100010 : data_out =  24'b000000001111111010010010;
		16'b0001011000100100 : data_out =  24'b000000001111111011010011;
		16'b0001011000100110 : data_out =  24'b000000001111111100010101;
		16'b0001011000101000 : data_out =  24'b000000001111111101010110;
		16'b0001011000101011 : data_out =  24'b000000001111111110010111;
		16'b0001011000101101 : data_out =  24'b000000001111111111011001;
		16'b0001011000101111 : data_out =  24'b000000010000000000011010;
		16'b0001011000110001 : data_out =  24'b000000010000000001011100;
		16'b0001011000110011 : data_out =  24'b000000010000000010011110;
		16'b0001011000110101 : data_out =  24'b000000010000000011011111;
		16'b0001011000110111 : data_out =  24'b000000010000000100100001;
		16'b0001011000111001 : data_out =  24'b000000010000000101100011;
		16'b0001011000111011 : data_out =  24'b000000010000000110100101;
		16'b0001011000111101 : data_out =  24'b000000010000000111100111;
		16'b0001011000111111 : data_out =  24'b000000010000001000101001;
		16'b0001011001000001 : data_out =  24'b000000010000001001101011;
		16'b0001011001000011 : data_out =  24'b000000010000001010101101;
		16'b0001011001000101 : data_out =  24'b000000010000001011110000;
		16'b0001011001000111 : data_out =  24'b000000010000001100110010;
		16'b0001011001001001 : data_out =  24'b000000010000001101110100;
		16'b0001011001001011 : data_out =  24'b000000010000001110110111;
		16'b0001011001001101 : data_out =  24'b000000010000001111111001;
		16'b0001011001001111 : data_out =  24'b000000010000010000111100;
		16'b0001011001010001 : data_out =  24'b000000010000010001111111;
		16'b0001011001010011 : data_out =  24'b000000010000010011000001;
		16'b0001011001010110 : data_out =  24'b000000010000010100000100;
		16'b0001011001011000 : data_out =  24'b000000010000010101000111;
		16'b0001011001011010 : data_out =  24'b000000010000010110001010;
		16'b0001011001011100 : data_out =  24'b000000010000010111001101;
		16'b0001011001011110 : data_out =  24'b000000010000011000010000;
		16'b0001011001100000 : data_out =  24'b000000010000011001010011;
		16'b0001011001100010 : data_out =  24'b000000010000011010010110;
		16'b0001011001100100 : data_out =  24'b000000010000011011011001;
		16'b0001011001100110 : data_out =  24'b000000010000011100011101;
		16'b0001011001101000 : data_out =  24'b000000010000011101100000;
		16'b0001011001101010 : data_out =  24'b000000010000011110100100;
		16'b0001011001101100 : data_out =  24'b000000010000011111100111;
		16'b0001011001101110 : data_out =  24'b000000010000100000101011;
		16'b0001011001110000 : data_out =  24'b000000010000100001101110;
		16'b0001011001110010 : data_out =  24'b000000010000100010110010;
		16'b0001011001110100 : data_out =  24'b000000010000100011110110;
		16'b0001011001110110 : data_out =  24'b000000010000100100111010;
		16'b0001011001111000 : data_out =  24'b000000010000100101111110;
		16'b0001011001111010 : data_out =  24'b000000010000100111000010;
		16'b0001011001111100 : data_out =  24'b000000010000101000000110;
		16'b0001011001111110 : data_out =  24'b000000010000101001001010;
		16'b0001011010000001 : data_out =  24'b000000010000101010001110;
		16'b0001011010000011 : data_out =  24'b000000010000101011010010;
		16'b0001011010000101 : data_out =  24'b000000010000101100010111;
		16'b0001011010000111 : data_out =  24'b000000010000101101011011;
		16'b0001011010001001 : data_out =  24'b000000010000101110100000;
		16'b0001011010001011 : data_out =  24'b000000010000101111100100;
		16'b0001011010001101 : data_out =  24'b000000010000110000101001;
		16'b0001011010001111 : data_out =  24'b000000010000110001101101;
		16'b0001011010010001 : data_out =  24'b000000010000110010110010;
		16'b0001011010010011 : data_out =  24'b000000010000110011110111;
		16'b0001011010010101 : data_out =  24'b000000010000110100111100;
		16'b0001011010010111 : data_out =  24'b000000010000110110000001;
		16'b0001011010011001 : data_out =  24'b000000010000110111000110;
		16'b0001011010011011 : data_out =  24'b000000010000111000001011;
		16'b0001011010011101 : data_out =  24'b000000010000111001010000;
		16'b0001011010011111 : data_out =  24'b000000010000111010010101;
		16'b0001011010100001 : data_out =  24'b000000010000111011011011;
		16'b0001011010100011 : data_out =  24'b000000010000111100100000;
		16'b0001011010100101 : data_out =  24'b000000010000111101100110;
		16'b0001011010100111 : data_out =  24'b000000010000111110101011;
		16'b0001011010101001 : data_out =  24'b000000010000111111110001;
		16'b0001011010101100 : data_out =  24'b000000010001000000110110;
		16'b0001011010101110 : data_out =  24'b000000010001000001111100;
		16'b0001011010110000 : data_out =  24'b000000010001000011000010;
		16'b0001011010110010 : data_out =  24'b000000010001000100001000;
		16'b0001011010110100 : data_out =  24'b000000010001000101001110;
		16'b0001011010110110 : data_out =  24'b000000010001000110010100;
		16'b0001011010111000 : data_out =  24'b000000010001000111011010;
		16'b0001011010111010 : data_out =  24'b000000010001001000100000;
		16'b0001011010111100 : data_out =  24'b000000010001001001100110;
		16'b0001011010111110 : data_out =  24'b000000010001001010101100;
		16'b0001011011000000 : data_out =  24'b000000010001001011110011;
		16'b0001011011000010 : data_out =  24'b000000010001001100111001;
		16'b0001011011000100 : data_out =  24'b000000010001001110000000;
		16'b0001011011000110 : data_out =  24'b000000010001001111000110;
		16'b0001011011001000 : data_out =  24'b000000010001010000001101;
		16'b0001011011001010 : data_out =  24'b000000010001010001010011;
		16'b0001011011001100 : data_out =  24'b000000010001010010011010;
		16'b0001011011001110 : data_out =  24'b000000010001010011100001;
		16'b0001011011010000 : data_out =  24'b000000010001010100101000;
		16'b0001011011010010 : data_out =  24'b000000010001010101101111;
		16'b0001011011010100 : data_out =  24'b000000010001010110110110;
		16'b0001011011010111 : data_out =  24'b000000010001010111111101;
		16'b0001011011011001 : data_out =  24'b000000010001011001000100;
		16'b0001011011011011 : data_out =  24'b000000010001011010001100;
		16'b0001011011011101 : data_out =  24'b000000010001011011010011;
		16'b0001011011011111 : data_out =  24'b000000010001011100011010;
		16'b0001011011100001 : data_out =  24'b000000010001011101100010;
		16'b0001011011100011 : data_out =  24'b000000010001011110101001;
		16'b0001011011100101 : data_out =  24'b000000010001011111110001;
		16'b0001011011100111 : data_out =  24'b000000010001100000111001;
		16'b0001011011101001 : data_out =  24'b000000010001100010000001;
		16'b0001011011101011 : data_out =  24'b000000010001100011001000;
		16'b0001011011101101 : data_out =  24'b000000010001100100010000;
		16'b0001011011101111 : data_out =  24'b000000010001100101011000;
		16'b0001011011110001 : data_out =  24'b000000010001100110100000;
		16'b0001011011110011 : data_out =  24'b000000010001100111101001;
		16'b0001011011110101 : data_out =  24'b000000010001101000110001;
		16'b0001011011110111 : data_out =  24'b000000010001101001111001;
		16'b0001011011111001 : data_out =  24'b000000010001101011000001;
		16'b0001011011111011 : data_out =  24'b000000010001101100001010;
		16'b0001011011111101 : data_out =  24'b000000010001101101010010;
		16'b0001011011111111 : data_out =  24'b000000010001101110011011;
		16'b0001011100000010 : data_out =  24'b000000010001101111100011;
		16'b0001011100000100 : data_out =  24'b000000010001110000101100;
		16'b0001011100000110 : data_out =  24'b000000010001110001110101;
		16'b0001011100001000 : data_out =  24'b000000010001110010111110;
		16'b0001011100001010 : data_out =  24'b000000010001110100000111;
		16'b0001011100001100 : data_out =  24'b000000010001110101010000;
		16'b0001011100001110 : data_out =  24'b000000010001110110011001;
		16'b0001011100010000 : data_out =  24'b000000010001110111100010;
		16'b0001011100010010 : data_out =  24'b000000010001111000101011;
		16'b0001011100010100 : data_out =  24'b000000010001111001110101;
		16'b0001011100010110 : data_out =  24'b000000010001111010111110;
		16'b0001011100011000 : data_out =  24'b000000010001111100000111;
		16'b0001011100011010 : data_out =  24'b000000010001111101010001;
		16'b0001011100011100 : data_out =  24'b000000010001111110011010;
		16'b0001011100011110 : data_out =  24'b000000010001111111100100;
		16'b0001011100100000 : data_out =  24'b000000010010000000101110;
		16'b0001011100100010 : data_out =  24'b000000010010000001111000;
		16'b0001011100100100 : data_out =  24'b000000010010000011000010;
		16'b0001011100100110 : data_out =  24'b000000010010000100001011;
		16'b0001011100101000 : data_out =  24'b000000010010000101010110;
		16'b0001011100101011 : data_out =  24'b000000010010000110100000;
		16'b0001011100101101 : data_out =  24'b000000010010000111101010;
		16'b0001011100101111 : data_out =  24'b000000010010001000110100;
		16'b0001011100110001 : data_out =  24'b000000010010001001111110;
		16'b0001011100110011 : data_out =  24'b000000010010001011001001;
		16'b0001011100110101 : data_out =  24'b000000010010001100010011;
		16'b0001011100110111 : data_out =  24'b000000010010001101011110;
		16'b0001011100111001 : data_out =  24'b000000010010001110101000;
		16'b0001011100111011 : data_out =  24'b000000010010001111110011;
		16'b0001011100111101 : data_out =  24'b000000010010010000111110;
		16'b0001011100111111 : data_out =  24'b000000010010010010001001;
		16'b0001011101000001 : data_out =  24'b000000010010010011010100;
		16'b0001011101000011 : data_out =  24'b000000010010010100011111;
		16'b0001011101000101 : data_out =  24'b000000010010010101101010;
		16'b0001011101000111 : data_out =  24'b000000010010010110110101;
		16'b0001011101001001 : data_out =  24'b000000010010011000000000;
		16'b0001011101001011 : data_out =  24'b000000010010011001001011;
		16'b0001011101001101 : data_out =  24'b000000010010011010010111;
		16'b0001011101001111 : data_out =  24'b000000010010011011100010;
		16'b0001011101010001 : data_out =  24'b000000010010011100101110;
		16'b0001011101010011 : data_out =  24'b000000010010011101111001;
		16'b0001011101010110 : data_out =  24'b000000010010011111000101;
		16'b0001011101011000 : data_out =  24'b000000010010100000010001;
		16'b0001011101011010 : data_out =  24'b000000010010100001011101;
		16'b0001011101011100 : data_out =  24'b000000010010100010101001;
		16'b0001011101011110 : data_out =  24'b000000010010100011110101;
		16'b0001011101100000 : data_out =  24'b000000010010100101000001;
		16'b0001011101100010 : data_out =  24'b000000010010100110001101;
		16'b0001011101100100 : data_out =  24'b000000010010100111011001;
		16'b0001011101100110 : data_out =  24'b000000010010101000100101;
		16'b0001011101101000 : data_out =  24'b000000010010101001110010;
		16'b0001011101101010 : data_out =  24'b000000010010101010111110;
		16'b0001011101101100 : data_out =  24'b000000010010101100001011;
		16'b0001011101101110 : data_out =  24'b000000010010101101010111;
		16'b0001011101110000 : data_out =  24'b000000010010101110100100;
		16'b0001011101110010 : data_out =  24'b000000010010101111110001;
		16'b0001011101110100 : data_out =  24'b000000010010110000111101;
		16'b0001011101110110 : data_out =  24'b000000010010110010001010;
		16'b0001011101111000 : data_out =  24'b000000010010110011010111;
		16'b0001011101111010 : data_out =  24'b000000010010110100100100;
		16'b0001011101111100 : data_out =  24'b000000010010110101110010;
		16'b0001011101111110 : data_out =  24'b000000010010110110111111;
		16'b0001011110000001 : data_out =  24'b000000010010111000001100;
		16'b0001011110000011 : data_out =  24'b000000010010111001011001;
		16'b0001011110000101 : data_out =  24'b000000010010111010100111;
		16'b0001011110000111 : data_out =  24'b000000010010111011110100;
		16'b0001011110001001 : data_out =  24'b000000010010111101000010;
		16'b0001011110001011 : data_out =  24'b000000010010111110010000;
		16'b0001011110001101 : data_out =  24'b000000010010111111011101;
		16'b0001011110001111 : data_out =  24'b000000010011000000101011;
		16'b0001011110010001 : data_out =  24'b000000010011000001111001;
		16'b0001011110010011 : data_out =  24'b000000010011000011000111;
		16'b0001011110010101 : data_out =  24'b000000010011000100010101;
		16'b0001011110010111 : data_out =  24'b000000010011000101100011;
		16'b0001011110011001 : data_out =  24'b000000010011000110110001;
		16'b0001011110011011 : data_out =  24'b000000010011001000000000;
		16'b0001011110011101 : data_out =  24'b000000010011001001001110;
		16'b0001011110011111 : data_out =  24'b000000010011001010011101;
		16'b0001011110100001 : data_out =  24'b000000010011001011101011;
		16'b0001011110100011 : data_out =  24'b000000010011001100111010;
		16'b0001011110100101 : data_out =  24'b000000010011001110001000;
		16'b0001011110100111 : data_out =  24'b000000010011001111010111;
		16'b0001011110101001 : data_out =  24'b000000010011010000100110;
		16'b0001011110101100 : data_out =  24'b000000010011010001110101;
		16'b0001011110101110 : data_out =  24'b000000010011010011000100;
		16'b0001011110110000 : data_out =  24'b000000010011010100010011;
		16'b0001011110110010 : data_out =  24'b000000010011010101100010;
		16'b0001011110110100 : data_out =  24'b000000010011010110110001;
		16'b0001011110110110 : data_out =  24'b000000010011011000000001;
		16'b0001011110111000 : data_out =  24'b000000010011011001010000;
		16'b0001011110111010 : data_out =  24'b000000010011011010100000;
		16'b0001011110111100 : data_out =  24'b000000010011011011101111;
		16'b0001011110111110 : data_out =  24'b000000010011011100111111;
		16'b0001011111000000 : data_out =  24'b000000010011011110001111;
		16'b0001011111000010 : data_out =  24'b000000010011011111011110;
		16'b0001011111000100 : data_out =  24'b000000010011100000101110;
		16'b0001011111000110 : data_out =  24'b000000010011100001111110;
		16'b0001011111001000 : data_out =  24'b000000010011100011001110;
		16'b0001011111001010 : data_out =  24'b000000010011100100011110;
		16'b0001011111001100 : data_out =  24'b000000010011100101101111;
		16'b0001011111001110 : data_out =  24'b000000010011100110111111;
		16'b0001011111010000 : data_out =  24'b000000010011101000001111;
		16'b0001011111010010 : data_out =  24'b000000010011101001100000;
		16'b0001011111010100 : data_out =  24'b000000010011101010110000;
		16'b0001011111010111 : data_out =  24'b000000010011101100000001;
		16'b0001011111011001 : data_out =  24'b000000010011101101010001;
		16'b0001011111011011 : data_out =  24'b000000010011101110100010;
		16'b0001011111011101 : data_out =  24'b000000010011101111110011;
		16'b0001011111011111 : data_out =  24'b000000010011110001000100;
		16'b0001011111100001 : data_out =  24'b000000010011110010010101;
		16'b0001011111100011 : data_out =  24'b000000010011110011100110;
		16'b0001011111100101 : data_out =  24'b000000010011110100110111;
		16'b0001011111100111 : data_out =  24'b000000010011110110001001;
		16'b0001011111101001 : data_out =  24'b000000010011110111011010;
		16'b0001011111101011 : data_out =  24'b000000010011111000101011;
		16'b0001011111101101 : data_out =  24'b000000010011111001111101;
		16'b0001011111101111 : data_out =  24'b000000010011111011001110;
		16'b0001011111110001 : data_out =  24'b000000010011111100100000;
		16'b0001011111110011 : data_out =  24'b000000010011111101110010;
		16'b0001011111110101 : data_out =  24'b000000010011111111000100;
		16'b0001011111110111 : data_out =  24'b000000010100000000010101;
		16'b0001011111111001 : data_out =  24'b000000010100000001100111;
		16'b0001011111111011 : data_out =  24'b000000010100000010111001;
		16'b0001011111111101 : data_out =  24'b000000010100000100001100;
		16'b0001011111111111 : data_out =  24'b000000010100000101011110;
		16'b0001100000000010 : data_out =  24'b000000010100000110110000;
		16'b0001100000000100 : data_out =  24'b000000010100001000000011;
		16'b0001100000000110 : data_out =  24'b000000010100001001010101;
		16'b0001100000001000 : data_out =  24'b000000010100001010101000;
		16'b0001100000001010 : data_out =  24'b000000010100001011111010;
		16'b0001100000001100 : data_out =  24'b000000010100001101001101;
		16'b0001100000001110 : data_out =  24'b000000010100001110100000;
		16'b0001100000010000 : data_out =  24'b000000010100001111110011;
		16'b0001100000010010 : data_out =  24'b000000010100010001000110;
		16'b0001100000010100 : data_out =  24'b000000010100010010011001;
		16'b0001100000010110 : data_out =  24'b000000010100010011101100;
		16'b0001100000011000 : data_out =  24'b000000010100010100111111;
		16'b0001100000011010 : data_out =  24'b000000010100010110010010;
		16'b0001100000011100 : data_out =  24'b000000010100010111100110;
		16'b0001100000011110 : data_out =  24'b000000010100011000111001;
		16'b0001100000100000 : data_out =  24'b000000010100011010001101;
		16'b0001100000100010 : data_out =  24'b000000010100011011100000;
		16'b0001100000100100 : data_out =  24'b000000010100011100110100;
		16'b0001100000100110 : data_out =  24'b000000010100011110001000;
		16'b0001100000101000 : data_out =  24'b000000010100011111011100;
		16'b0001100000101011 : data_out =  24'b000000010100100000110000;
		16'b0001100000101101 : data_out =  24'b000000010100100010000100;
		16'b0001100000101111 : data_out =  24'b000000010100100011011000;
		16'b0001100000110001 : data_out =  24'b000000010100100100101100;
		16'b0001100000110011 : data_out =  24'b000000010100100110000001;
		16'b0001100000110101 : data_out =  24'b000000010100100111010101;
		16'b0001100000110111 : data_out =  24'b000000010100101000101001;
		16'b0001100000111001 : data_out =  24'b000000010100101001111110;
		16'b0001100000111011 : data_out =  24'b000000010100101011010011;
		16'b0001100000111101 : data_out =  24'b000000010100101100100111;
		16'b0001100000111111 : data_out =  24'b000000010100101101111100;
		16'b0001100001000001 : data_out =  24'b000000010100101111010001;
		16'b0001100001000011 : data_out =  24'b000000010100110000100110;
		16'b0001100001000101 : data_out =  24'b000000010100110001111011;
		16'b0001100001000111 : data_out =  24'b000000010100110011010000;
		16'b0001100001001001 : data_out =  24'b000000010100110100100110;
		16'b0001100001001011 : data_out =  24'b000000010100110101111011;
		16'b0001100001001101 : data_out =  24'b000000010100110111010000;
		16'b0001100001001111 : data_out =  24'b000000010100111000100110;
		16'b0001100001010001 : data_out =  24'b000000010100111001111011;
		16'b0001100001010011 : data_out =  24'b000000010100111011010001;
		16'b0001100001010110 : data_out =  24'b000000010100111100100111;
		16'b0001100001011000 : data_out =  24'b000000010100111101111101;
		16'b0001100001011010 : data_out =  24'b000000010100111111010011;
		16'b0001100001011100 : data_out =  24'b000000010101000000101001;
		16'b0001100001011110 : data_out =  24'b000000010101000001111111;
		16'b0001100001100000 : data_out =  24'b000000010101000011010101;
		16'b0001100001100010 : data_out =  24'b000000010101000100101011;
		16'b0001100001100100 : data_out =  24'b000000010101000110000010;
		16'b0001100001100110 : data_out =  24'b000000010101000111011000;
		16'b0001100001101000 : data_out =  24'b000000010101001000101110;
		16'b0001100001101010 : data_out =  24'b000000010101001010000101;
		16'b0001100001101100 : data_out =  24'b000000010101001011011100;
		16'b0001100001101110 : data_out =  24'b000000010101001100110011;
		16'b0001100001110000 : data_out =  24'b000000010101001110001001;
		16'b0001100001110010 : data_out =  24'b000000010101001111100000;
		16'b0001100001110100 : data_out =  24'b000000010101010000110111;
		16'b0001100001110110 : data_out =  24'b000000010101010010001111;
		16'b0001100001111000 : data_out =  24'b000000010101010011100110;
		16'b0001100001111010 : data_out =  24'b000000010101010100111101;
		16'b0001100001111100 : data_out =  24'b000000010101010110010101;
		16'b0001100001111110 : data_out =  24'b000000010101010111101100;
		16'b0001100010000001 : data_out =  24'b000000010101011001000100;
		16'b0001100010000011 : data_out =  24'b000000010101011010011011;
		16'b0001100010000101 : data_out =  24'b000000010101011011110011;
		16'b0001100010000111 : data_out =  24'b000000010101011101001011;
		16'b0001100010001001 : data_out =  24'b000000010101011110100011;
		16'b0001100010001011 : data_out =  24'b000000010101011111111011;
		16'b0001100010001101 : data_out =  24'b000000010101100001010011;
		16'b0001100010001111 : data_out =  24'b000000010101100010101011;
		16'b0001100010010001 : data_out =  24'b000000010101100100000011;
		16'b0001100010010011 : data_out =  24'b000000010101100101011100;
		16'b0001100010010101 : data_out =  24'b000000010101100110110100;
		16'b0001100010010111 : data_out =  24'b000000010101101000001101;
		16'b0001100010011001 : data_out =  24'b000000010101101001100101;
		16'b0001100010011011 : data_out =  24'b000000010101101010111110;
		16'b0001100010011101 : data_out =  24'b000000010101101100010111;
		16'b0001100010011111 : data_out =  24'b000000010101101101110000;
		16'b0001100010100001 : data_out =  24'b000000010101101111001001;
		16'b0001100010100011 : data_out =  24'b000000010101110000100010;
		16'b0001100010100101 : data_out =  24'b000000010101110001111011;
		16'b0001100010100111 : data_out =  24'b000000010101110011010100;
		16'b0001100010101001 : data_out =  24'b000000010101110100101110;
		16'b0001100010101100 : data_out =  24'b000000010101110110000111;
		16'b0001100010101110 : data_out =  24'b000000010101110111100001;
		16'b0001100010110000 : data_out =  24'b000000010101111000111010;
		16'b0001100010110010 : data_out =  24'b000000010101111010010100;
		16'b0001100010110100 : data_out =  24'b000000010101111011101110;
		16'b0001100010110110 : data_out =  24'b000000010101111101001000;
		16'b0001100010111000 : data_out =  24'b000000010101111110100010;
		16'b0001100010111010 : data_out =  24'b000000010101111111111100;
		16'b0001100010111100 : data_out =  24'b000000010110000001010110;
		16'b0001100010111110 : data_out =  24'b000000010110000010110000;
		16'b0001100011000000 : data_out =  24'b000000010110000100001010;
		16'b0001100011000010 : data_out =  24'b000000010110000101100101;
		16'b0001100011000100 : data_out =  24'b000000010110000110111111;
		16'b0001100011000110 : data_out =  24'b000000010110001000011010;
		16'b0001100011001000 : data_out =  24'b000000010110001001110101;
		16'b0001100011001010 : data_out =  24'b000000010110001011001111;
		16'b0001100011001100 : data_out =  24'b000000010110001100101010;
		16'b0001100011001110 : data_out =  24'b000000010110001110000101;
		16'b0001100011010000 : data_out =  24'b000000010110001111100000;
		16'b0001100011010010 : data_out =  24'b000000010110010000111011;
		16'b0001100011010100 : data_out =  24'b000000010110010010010111;
		16'b0001100011010111 : data_out =  24'b000000010110010011110010;
		16'b0001100011011001 : data_out =  24'b000000010110010101001101;
		16'b0001100011011011 : data_out =  24'b000000010110010110101001;
		16'b0001100011011101 : data_out =  24'b000000010110011000000101;
		16'b0001100011011111 : data_out =  24'b000000010110011001100000;
		16'b0001100011100001 : data_out =  24'b000000010110011010111100;
		16'b0001100011100011 : data_out =  24'b000000010110011100011000;
		16'b0001100011100101 : data_out =  24'b000000010110011101110100;
		16'b0001100011100111 : data_out =  24'b000000010110011111010000;
		16'b0001100011101001 : data_out =  24'b000000010110100000101100;
		16'b0001100011101011 : data_out =  24'b000000010110100010001000;
		16'b0001100011101101 : data_out =  24'b000000010110100011100101;
		16'b0001100011101111 : data_out =  24'b000000010110100101000001;
		16'b0001100011110001 : data_out =  24'b000000010110100110011110;
		16'b0001100011110011 : data_out =  24'b000000010110100111111010;
		16'b0001100011110101 : data_out =  24'b000000010110101001010111;
		16'b0001100011110111 : data_out =  24'b000000010110101010110100;
		16'b0001100011111001 : data_out =  24'b000000010110101100010001;
		16'b0001100011111011 : data_out =  24'b000000010110101101101110;
		16'b0001100011111101 : data_out =  24'b000000010110101111001011;
		16'b0001100011111111 : data_out =  24'b000000010110110000101000;
		16'b0001100100000010 : data_out =  24'b000000010110110010000101;
		16'b0001100100000100 : data_out =  24'b000000010110110011100011;
		16'b0001100100000110 : data_out =  24'b000000010110110101000000;
		16'b0001100100001000 : data_out =  24'b000000010110110110011110;
		16'b0001100100001010 : data_out =  24'b000000010110110111111011;
		16'b0001100100001100 : data_out =  24'b000000010110111001011001;
		16'b0001100100001110 : data_out =  24'b000000010110111010110111;
		16'b0001100100010000 : data_out =  24'b000000010110111100010101;
		16'b0001100100010010 : data_out =  24'b000000010110111101110011;
		16'b0001100100010100 : data_out =  24'b000000010110111111010001;
		16'b0001100100010110 : data_out =  24'b000000010111000000101111;
		16'b0001100100011000 : data_out =  24'b000000010111000010001101;
		16'b0001100100011010 : data_out =  24'b000000010111000011101100;
		16'b0001100100011100 : data_out =  24'b000000010111000101001010;
		16'b0001100100011110 : data_out =  24'b000000010111000110101001;
		16'b0001100100100000 : data_out =  24'b000000010111001000001000;
		16'b0001100100100010 : data_out =  24'b000000010111001001100110;
		16'b0001100100100100 : data_out =  24'b000000010111001011000101;
		16'b0001100100100110 : data_out =  24'b000000010111001100100100;
		16'b0001100100101000 : data_out =  24'b000000010111001110000011;
		16'b0001100100101011 : data_out =  24'b000000010111001111100010;
		16'b0001100100101101 : data_out =  24'b000000010111010001000010;
		16'b0001100100101111 : data_out =  24'b000000010111010010100001;
		16'b0001100100110001 : data_out =  24'b000000010111010100000000;
		16'b0001100100110011 : data_out =  24'b000000010111010101100000;
		16'b0001100100110101 : data_out =  24'b000000010111010111000000;
		16'b0001100100110111 : data_out =  24'b000000010111011000011111;
		16'b0001100100111001 : data_out =  24'b000000010111011001111111;
		16'b0001100100111011 : data_out =  24'b000000010111011011011111;
		16'b0001100100111101 : data_out =  24'b000000010111011100111111;
		16'b0001100100111111 : data_out =  24'b000000010111011110011111;
		16'b0001100101000001 : data_out =  24'b000000010111011111111111;
		16'b0001100101000011 : data_out =  24'b000000010111100001100000;
		16'b0001100101000101 : data_out =  24'b000000010111100011000000;
		16'b0001100101000111 : data_out =  24'b000000010111100100100001;
		16'b0001100101001001 : data_out =  24'b000000010111100110000001;
		16'b0001100101001011 : data_out =  24'b000000010111100111100010;
		16'b0001100101001101 : data_out =  24'b000000010111101001000011;
		16'b0001100101001111 : data_out =  24'b000000010111101010100100;
		16'b0001100101010001 : data_out =  24'b000000010111101100000101;
		16'b0001100101010011 : data_out =  24'b000000010111101101100110;
		16'b0001100101010110 : data_out =  24'b000000010111101111000111;
		16'b0001100101011000 : data_out =  24'b000000010111110000101000;
		16'b0001100101011010 : data_out =  24'b000000010111110010001001;
		16'b0001100101011100 : data_out =  24'b000000010111110011101011;
		16'b0001100101011110 : data_out =  24'b000000010111110101001101;
		16'b0001100101100000 : data_out =  24'b000000010111110110101110;
		16'b0001100101100010 : data_out =  24'b000000010111111000010000;
		16'b0001100101100100 : data_out =  24'b000000010111111001110010;
		16'b0001100101100110 : data_out =  24'b000000010111111011010100;
		16'b0001100101101000 : data_out =  24'b000000010111111100110110;
		16'b0001100101101010 : data_out =  24'b000000010111111110011000;
		16'b0001100101101100 : data_out =  24'b000000010111111111111010;
		16'b0001100101101110 : data_out =  24'b000000011000000001011101;
		16'b0001100101110000 : data_out =  24'b000000011000000010111111;
		16'b0001100101110010 : data_out =  24'b000000011000000100100010;
		16'b0001100101110100 : data_out =  24'b000000011000000110000100;
		16'b0001100101110110 : data_out =  24'b000000011000000111100111;
		16'b0001100101111000 : data_out =  24'b000000011000001001001010;
		16'b0001100101111010 : data_out =  24'b000000011000001010101101;
		16'b0001100101111100 : data_out =  24'b000000011000001100010000;
		16'b0001100101111110 : data_out =  24'b000000011000001101110011;
		16'b0001100110000001 : data_out =  24'b000000011000001111010110;
		16'b0001100110000011 : data_out =  24'b000000011000010000111001;
		16'b0001100110000101 : data_out =  24'b000000011000010010011101;
		16'b0001100110000111 : data_out =  24'b000000011000010100000000;
		16'b0001100110001001 : data_out =  24'b000000011000010101100100;
		16'b0001100110001011 : data_out =  24'b000000011000010111001000;
		16'b0001100110001101 : data_out =  24'b000000011000011000101100;
		16'b0001100110001111 : data_out =  24'b000000011000011010010000;
		16'b0001100110010001 : data_out =  24'b000000011000011011110100;
		16'b0001100110010011 : data_out =  24'b000000011000011101011000;
		16'b0001100110010101 : data_out =  24'b000000011000011110111100;
		16'b0001100110010111 : data_out =  24'b000000011000100000100000;
		16'b0001100110011001 : data_out =  24'b000000011000100010000101;
		16'b0001100110011011 : data_out =  24'b000000011000100011101001;
		16'b0001100110011101 : data_out =  24'b000000011000100101001110;
		16'b0001100110011111 : data_out =  24'b000000011000100110110011;
		16'b0001100110100001 : data_out =  24'b000000011000101000010111;
		16'b0001100110100011 : data_out =  24'b000000011000101001111100;
		16'b0001100110100101 : data_out =  24'b000000011000101011100001;
		16'b0001100110100111 : data_out =  24'b000000011000101101000111;
		16'b0001100110101001 : data_out =  24'b000000011000101110101100;
		16'b0001100110101100 : data_out =  24'b000000011000110000010001;
		16'b0001100110101110 : data_out =  24'b000000011000110001110111;
		16'b0001100110110000 : data_out =  24'b000000011000110011011100;
		16'b0001100110110010 : data_out =  24'b000000011000110101000010;
		16'b0001100110110100 : data_out =  24'b000000011000110110101000;
		16'b0001100110110110 : data_out =  24'b000000011000111000001101;
		16'b0001100110111000 : data_out =  24'b000000011000111001110011;
		16'b0001100110111010 : data_out =  24'b000000011000111011011001;
		16'b0001100110111100 : data_out =  24'b000000011000111101000000;
		16'b0001100110111110 : data_out =  24'b000000011000111110100110;
		16'b0001100111000000 : data_out =  24'b000000011001000000001100;
		16'b0001100111000010 : data_out =  24'b000000011001000001110011;
		16'b0001100111000100 : data_out =  24'b000000011001000011011001;
		16'b0001100111000110 : data_out =  24'b000000011001000101000000;
		16'b0001100111001000 : data_out =  24'b000000011001000110100111;
		16'b0001100111001010 : data_out =  24'b000000011001001000001110;
		16'b0001100111001100 : data_out =  24'b000000011001001001110101;
		16'b0001100111001110 : data_out =  24'b000000011001001011011100;
		16'b0001100111010000 : data_out =  24'b000000011001001101000011;
		16'b0001100111010010 : data_out =  24'b000000011001001110101010;
		16'b0001100111010100 : data_out =  24'b000000011001010000010001;
		16'b0001100111010111 : data_out =  24'b000000011001010001111001;
		16'b0001100111011001 : data_out =  24'b000000011001010011100001;
		16'b0001100111011011 : data_out =  24'b000000011001010101001000;
		16'b0001100111011101 : data_out =  24'b000000011001010110110000;
		16'b0001100111011111 : data_out =  24'b000000011001011000011000;
		16'b0001100111100001 : data_out =  24'b000000011001011010000000;
		16'b0001100111100011 : data_out =  24'b000000011001011011101000;
		16'b0001100111100101 : data_out =  24'b000000011001011101010000;
		16'b0001100111100111 : data_out =  24'b000000011001011110111001;
		16'b0001100111101001 : data_out =  24'b000000011001100000100001;
		16'b0001100111101011 : data_out =  24'b000000011001100010001010;
		16'b0001100111101101 : data_out =  24'b000000011001100011110010;
		16'b0001100111101111 : data_out =  24'b000000011001100101011011;
		16'b0001100111110001 : data_out =  24'b000000011001100111000100;
		16'b0001100111110011 : data_out =  24'b000000011001101000101101;
		16'b0001100111110101 : data_out =  24'b000000011001101010010110;
		16'b0001100111110111 : data_out =  24'b000000011001101011111111;
		16'b0001100111111001 : data_out =  24'b000000011001101101101000;
		16'b0001100111111011 : data_out =  24'b000000011001101111010010;
		16'b0001100111111101 : data_out =  24'b000000011001110000111011;
		16'b0001100111111111 : data_out =  24'b000000011001110010100101;
		16'b0001101000000010 : data_out =  24'b000000011001110100001110;
		16'b0001101000000100 : data_out =  24'b000000011001110101111000;
		16'b0001101000000110 : data_out =  24'b000000011001110111100010;
		16'b0001101000001000 : data_out =  24'b000000011001111001001100;
		16'b0001101000001010 : data_out =  24'b000000011001111010110110;
		16'b0001101000001100 : data_out =  24'b000000011001111100100000;
		16'b0001101000001110 : data_out =  24'b000000011001111110001011;
		16'b0001101000010000 : data_out =  24'b000000011001111111110101;
		16'b0001101000010010 : data_out =  24'b000000011010000001100000;
		16'b0001101000010100 : data_out =  24'b000000011010000011001010;
		16'b0001101000010110 : data_out =  24'b000000011010000100110101;
		16'b0001101000011000 : data_out =  24'b000000011010000110100000;
		16'b0001101000011010 : data_out =  24'b000000011010001000001011;
		16'b0001101000011100 : data_out =  24'b000000011010001001110110;
		16'b0001101000011110 : data_out =  24'b000000011010001011100001;
		16'b0001101000100000 : data_out =  24'b000000011010001101001101;
		16'b0001101000100010 : data_out =  24'b000000011010001110111000;
		16'b0001101000100100 : data_out =  24'b000000011010010000100011;
		16'b0001101000100110 : data_out =  24'b000000011010010010001111;
		16'b0001101000101000 : data_out =  24'b000000011010010011111011;
		16'b0001101000101011 : data_out =  24'b000000011010010101100111;
		16'b0001101000101101 : data_out =  24'b000000011010010111010011;
		16'b0001101000101111 : data_out =  24'b000000011010011000111111;
		16'b0001101000110001 : data_out =  24'b000000011010011010101011;
		16'b0001101000110011 : data_out =  24'b000000011010011100010111;
		16'b0001101000110101 : data_out =  24'b000000011010011110000011;
		16'b0001101000110111 : data_out =  24'b000000011010011111110000;
		16'b0001101000111001 : data_out =  24'b000000011010100001011100;
		16'b0001101000111011 : data_out =  24'b000000011010100011001001;
		16'b0001101000111101 : data_out =  24'b000000011010100100110110;
		16'b0001101000111111 : data_out =  24'b000000011010100110100011;
		16'b0001101001000001 : data_out =  24'b000000011010101000010000;
		16'b0001101001000011 : data_out =  24'b000000011010101001111101;
		16'b0001101001000101 : data_out =  24'b000000011010101011101010;
		16'b0001101001000111 : data_out =  24'b000000011010101101010111;
		16'b0001101001001001 : data_out =  24'b000000011010101111000101;
		16'b0001101001001011 : data_out =  24'b000000011010110000110011;
		16'b0001101001001101 : data_out =  24'b000000011010110010100000;
		16'b0001101001001111 : data_out =  24'b000000011010110100001110;
		16'b0001101001010001 : data_out =  24'b000000011010110101111100;
		16'b0001101001010011 : data_out =  24'b000000011010110111101010;
		16'b0001101001010110 : data_out =  24'b000000011010111001011000;
		16'b0001101001011000 : data_out =  24'b000000011010111011000110;
		16'b0001101001011010 : data_out =  24'b000000011010111100110101;
		16'b0001101001011100 : data_out =  24'b000000011010111110100011;
		16'b0001101001011110 : data_out =  24'b000000011011000000010010;
		16'b0001101001100000 : data_out =  24'b000000011011000010000000;
		16'b0001101001100010 : data_out =  24'b000000011011000011101111;
		16'b0001101001100100 : data_out =  24'b000000011011000101011110;
		16'b0001101001100110 : data_out =  24'b000000011011000111001101;
		16'b0001101001101000 : data_out =  24'b000000011011001000111100;
		16'b0001101001101010 : data_out =  24'b000000011011001010101011;
		16'b0001101001101100 : data_out =  24'b000000011011001100011011;
		16'b0001101001101110 : data_out =  24'b000000011011001110001010;
		16'b0001101001110000 : data_out =  24'b000000011011001111111010;
		16'b0001101001110010 : data_out =  24'b000000011011010001101001;
		16'b0001101001110100 : data_out =  24'b000000011011010011011001;
		16'b0001101001110110 : data_out =  24'b000000011011010101001001;
		16'b0001101001111000 : data_out =  24'b000000011011010110111001;
		16'b0001101001111010 : data_out =  24'b000000011011011000101001;
		16'b0001101001111100 : data_out =  24'b000000011011011010011001;
		16'b0001101001111110 : data_out =  24'b000000011011011100001010;
		16'b0001101010000001 : data_out =  24'b000000011011011101111010;
		16'b0001101010000011 : data_out =  24'b000000011011011111101011;
		16'b0001101010000101 : data_out =  24'b000000011011100001011011;
		16'b0001101010000111 : data_out =  24'b000000011011100011001100;
		16'b0001101010001001 : data_out =  24'b000000011011100100111101;
		16'b0001101010001011 : data_out =  24'b000000011011100110101110;
		16'b0001101010001101 : data_out =  24'b000000011011101000011111;
		16'b0001101010001111 : data_out =  24'b000000011011101010010000;
		16'b0001101010010001 : data_out =  24'b000000011011101100000010;
		16'b0001101010010011 : data_out =  24'b000000011011101101110011;
		16'b0001101010010101 : data_out =  24'b000000011011101111100101;
		16'b0001101010010111 : data_out =  24'b000000011011110001010110;
		16'b0001101010011001 : data_out =  24'b000000011011110011001000;
		16'b0001101010011011 : data_out =  24'b000000011011110100111010;
		16'b0001101010011101 : data_out =  24'b000000011011110110101100;
		16'b0001101010011111 : data_out =  24'b000000011011111000011110;
		16'b0001101010100001 : data_out =  24'b000000011011111010010001;
		16'b0001101010100011 : data_out =  24'b000000011011111100000011;
		16'b0001101010100101 : data_out =  24'b000000011011111101110101;
		16'b0001101010100111 : data_out =  24'b000000011011111111101000;
		16'b0001101010101001 : data_out =  24'b000000011100000001011011;
		16'b0001101010101100 : data_out =  24'b000000011100000011001110;
		16'b0001101010101110 : data_out =  24'b000000011100000101000001;
		16'b0001101010110000 : data_out =  24'b000000011100000110110100;
		16'b0001101010110010 : data_out =  24'b000000011100001000100111;
		16'b0001101010110100 : data_out =  24'b000000011100001010011010;
		16'b0001101010110110 : data_out =  24'b000000011100001100001110;
		16'b0001101010111000 : data_out =  24'b000000011100001110000001;
		16'b0001101010111010 : data_out =  24'b000000011100001111110101;
		16'b0001101010111100 : data_out =  24'b000000011100010001101000;
		16'b0001101010111110 : data_out =  24'b000000011100010011011100;
		16'b0001101011000000 : data_out =  24'b000000011100010101010000;
		16'b0001101011000010 : data_out =  24'b000000011100010111000100;
		16'b0001101011000100 : data_out =  24'b000000011100011000111001;
		16'b0001101011000110 : data_out =  24'b000000011100011010101101;
		16'b0001101011001000 : data_out =  24'b000000011100011100100001;
		16'b0001101011001010 : data_out =  24'b000000011100011110010110;
		16'b0001101011001100 : data_out =  24'b000000011100100000001011;
		16'b0001101011001110 : data_out =  24'b000000011100100010000000;
		16'b0001101011010000 : data_out =  24'b000000011100100011110100;
		16'b0001101011010010 : data_out =  24'b000000011100100101101001;
		16'b0001101011010100 : data_out =  24'b000000011100100111011111;
		16'b0001101011010111 : data_out =  24'b000000011100101001010100;
		16'b0001101011011001 : data_out =  24'b000000011100101011001001;
		16'b0001101011011011 : data_out =  24'b000000011100101100111111;
		16'b0001101011011101 : data_out =  24'b000000011100101110110100;
		16'b0001101011011111 : data_out =  24'b000000011100110000101010;
		16'b0001101011100001 : data_out =  24'b000000011100110010100000;
		16'b0001101011100011 : data_out =  24'b000000011100110100010110;
		16'b0001101011100101 : data_out =  24'b000000011100110110001100;
		16'b0001101011100111 : data_out =  24'b000000011100111000000010;
		16'b0001101011101001 : data_out =  24'b000000011100111001111001;
		16'b0001101011101011 : data_out =  24'b000000011100111011101111;
		16'b0001101011101101 : data_out =  24'b000000011100111101100110;
		16'b0001101011101111 : data_out =  24'b000000011100111111011100;
		16'b0001101011110001 : data_out =  24'b000000011101000001010011;
		16'b0001101011110011 : data_out =  24'b000000011101000011001010;
		16'b0001101011110101 : data_out =  24'b000000011101000101000001;
		16'b0001101011110111 : data_out =  24'b000000011101000110111000;
		16'b0001101011111001 : data_out =  24'b000000011101001000110000;
		16'b0001101011111011 : data_out =  24'b000000011101001010100111;
		16'b0001101011111101 : data_out =  24'b000000011101001100011111;
		16'b0001101011111111 : data_out =  24'b000000011101001110010110;
		16'b0001101100000010 : data_out =  24'b000000011101010000001110;
		16'b0001101100000100 : data_out =  24'b000000011101010010000110;
		16'b0001101100000110 : data_out =  24'b000000011101010011111110;
		16'b0001101100001000 : data_out =  24'b000000011101010101110110;
		16'b0001101100001010 : data_out =  24'b000000011101010111101110;
		16'b0001101100001100 : data_out =  24'b000000011101011001100111;
		16'b0001101100001110 : data_out =  24'b000000011101011011011111;
		16'b0001101100010000 : data_out =  24'b000000011101011101011000;
		16'b0001101100010010 : data_out =  24'b000000011101011111010000;
		16'b0001101100010100 : data_out =  24'b000000011101100001001001;
		16'b0001101100010110 : data_out =  24'b000000011101100011000010;
		16'b0001101100011000 : data_out =  24'b000000011101100100111011;
		16'b0001101100011010 : data_out =  24'b000000011101100110110100;
		16'b0001101100011100 : data_out =  24'b000000011101101000101110;
		16'b0001101100011110 : data_out =  24'b000000011101101010100111;
		16'b0001101100100000 : data_out =  24'b000000011101101100100001;
		16'b0001101100100010 : data_out =  24'b000000011101101110011011;
		16'b0001101100100100 : data_out =  24'b000000011101110000010100;
		16'b0001101100100110 : data_out =  24'b000000011101110010001110;
		16'b0001101100101000 : data_out =  24'b000000011101110100001000;
		16'b0001101100101011 : data_out =  24'b000000011101110110000011;
		16'b0001101100101101 : data_out =  24'b000000011101110111111101;
		16'b0001101100101111 : data_out =  24'b000000011101111001110111;
		16'b0001101100110001 : data_out =  24'b000000011101111011110010;
		16'b0001101100110011 : data_out =  24'b000000011101111101101100;
		16'b0001101100110101 : data_out =  24'b000000011101111111100111;
		16'b0001101100110111 : data_out =  24'b000000011110000001100010;
		16'b0001101100111001 : data_out =  24'b000000011110000011011101;
		16'b0001101100111011 : data_out =  24'b000000011110000101011000;
		16'b0001101100111101 : data_out =  24'b000000011110000111010100;
		16'b0001101100111111 : data_out =  24'b000000011110001001001111;
		16'b0001101101000001 : data_out =  24'b000000011110001011001011;
		16'b0001101101000011 : data_out =  24'b000000011110001101000110;
		16'b0001101101000101 : data_out =  24'b000000011110001111000010;
		16'b0001101101000111 : data_out =  24'b000000011110010000111110;
		16'b0001101101001001 : data_out =  24'b000000011110010010111010;
		16'b0001101101001011 : data_out =  24'b000000011110010100110110;
		16'b0001101101001101 : data_out =  24'b000000011110010110110010;
		16'b0001101101001111 : data_out =  24'b000000011110011000101111;
		16'b0001101101010001 : data_out =  24'b000000011110011010101011;
		16'b0001101101010011 : data_out =  24'b000000011110011100101000;
		16'b0001101101010110 : data_out =  24'b000000011110011110100101;
		16'b0001101101011000 : data_out =  24'b000000011110100000100010;
		16'b0001101101011010 : data_out =  24'b000000011110100010011111;
		16'b0001101101011100 : data_out =  24'b000000011110100100011100;
		16'b0001101101011110 : data_out =  24'b000000011110100110011001;
		16'b0001101101100000 : data_out =  24'b000000011110101000010110;
		16'b0001101101100010 : data_out =  24'b000000011110101010010100;
		16'b0001101101100100 : data_out =  24'b000000011110101100010010;
		16'b0001101101100110 : data_out =  24'b000000011110101110001111;
		16'b0001101101101000 : data_out =  24'b000000011110110000001101;
		16'b0001101101101010 : data_out =  24'b000000011110110010001011;
		16'b0001101101101100 : data_out =  24'b000000011110110100001010;
		16'b0001101101101110 : data_out =  24'b000000011110110110001000;
		16'b0001101101110000 : data_out =  24'b000000011110111000000110;
		16'b0001101101110010 : data_out =  24'b000000011110111010000101;
		16'b0001101101110100 : data_out =  24'b000000011110111100000011;
		16'b0001101101110110 : data_out =  24'b000000011110111110000010;
		16'b0001101101111000 : data_out =  24'b000000011111000000000001;
		16'b0001101101111010 : data_out =  24'b000000011111000010000000;
		16'b0001101101111100 : data_out =  24'b000000011111000011111111;
		16'b0001101101111110 : data_out =  24'b000000011111000101111111;
		16'b0001101110000001 : data_out =  24'b000000011111000111111110;
		16'b0001101110000011 : data_out =  24'b000000011111001001111110;
		16'b0001101110000101 : data_out =  24'b000000011111001011111101;
		16'b0001101110000111 : data_out =  24'b000000011111001101111101;
		16'b0001101110001001 : data_out =  24'b000000011111001111111101;
		16'b0001101110001011 : data_out =  24'b000000011111010001111101;
		16'b0001101110001101 : data_out =  24'b000000011111010011111101;
		16'b0001101110001111 : data_out =  24'b000000011111010101111110;
		16'b0001101110010001 : data_out =  24'b000000011111010111111110;
		16'b0001101110010011 : data_out =  24'b000000011111011001111111;
		16'b0001101110010101 : data_out =  24'b000000011111011011111111;
		16'b0001101110010111 : data_out =  24'b000000011111011110000000;
		16'b0001101110011001 : data_out =  24'b000000011111100000000001;
		16'b0001101110011011 : data_out =  24'b000000011111100010000010;
		16'b0001101110011101 : data_out =  24'b000000011111100100000011;
		16'b0001101110011111 : data_out =  24'b000000011111100110000101;
		16'b0001101110100001 : data_out =  24'b000000011111101000000110;
		16'b0001101110100011 : data_out =  24'b000000011111101010001000;
		16'b0001101110100101 : data_out =  24'b000000011111101100001010;
		16'b0001101110100111 : data_out =  24'b000000011111101110001011;
		16'b0001101110101001 : data_out =  24'b000000011111110000001101;
		16'b0001101110101100 : data_out =  24'b000000011111110010010000;
		16'b0001101110101110 : data_out =  24'b000000011111110100010010;
		16'b0001101110110000 : data_out =  24'b000000011111110110010100;
		16'b0001101110110010 : data_out =  24'b000000011111111000010111;
		16'b0001101110110100 : data_out =  24'b000000011111111010011001;
		16'b0001101110110110 : data_out =  24'b000000011111111100011100;
		16'b0001101110111000 : data_out =  24'b000000011111111110011111;
		16'b0001101110111010 : data_out =  24'b000000100000000000100010;
		16'b0001101110111100 : data_out =  24'b000000100000000010100101;
		16'b0001101110111110 : data_out =  24'b000000100000000100101001;
		16'b0001101111000000 : data_out =  24'b000000100000000110101100;
		16'b0001101111000010 : data_out =  24'b000000100000001000110000;
		16'b0001101111000100 : data_out =  24'b000000100000001010110011;
		16'b0001101111000110 : data_out =  24'b000000100000001100110111;
		16'b0001101111001000 : data_out =  24'b000000100000001110111011;
		16'b0001101111001010 : data_out =  24'b000000100000010000111111;
		16'b0001101111001100 : data_out =  24'b000000100000010011000011;
		16'b0001101111001110 : data_out =  24'b000000100000010101001000;
		16'b0001101111010000 : data_out =  24'b000000100000010111001100;
		16'b0001101111010010 : data_out =  24'b000000100000011001010001;
		16'b0001101111010100 : data_out =  24'b000000100000011011010110;
		16'b0001101111010111 : data_out =  24'b000000100000011101011011;
		16'b0001101111011001 : data_out =  24'b000000100000011111100000;
		16'b0001101111011011 : data_out =  24'b000000100000100001100101;
		16'b0001101111011101 : data_out =  24'b000000100000100011101010;
		16'b0001101111011111 : data_out =  24'b000000100000100101101111;
		16'b0001101111100001 : data_out =  24'b000000100000100111110101;
		16'b0001101111100011 : data_out =  24'b000000100000101001111011;
		16'b0001101111100101 : data_out =  24'b000000100000101100000000;
		16'b0001101111100111 : data_out =  24'b000000100000101110000110;
		16'b0001101111101001 : data_out =  24'b000000100000110000001101;
		16'b0001101111101011 : data_out =  24'b000000100000110010010011;
		16'b0001101111101101 : data_out =  24'b000000100000110100011001;
		16'b0001101111101111 : data_out =  24'b000000100000110110100000;
		16'b0001101111110001 : data_out =  24'b000000100000111000100110;
		16'b0001101111110011 : data_out =  24'b000000100000111010101101;
		16'b0001101111110101 : data_out =  24'b000000100000111100110100;
		16'b0001101111110111 : data_out =  24'b000000100000111110111011;
		16'b0001101111111001 : data_out =  24'b000000100001000001000010;
		16'b0001101111111011 : data_out =  24'b000000100001000011001001;
		16'b0001101111111101 : data_out =  24'b000000100001000101010001;
		16'b0001101111111111 : data_out =  24'b000000100001000111011000;
		16'b0001110000000010 : data_out =  24'b000000100001001001100000;
		16'b0001110000000100 : data_out =  24'b000000100001001011101000;
		16'b0001110000000110 : data_out =  24'b000000100001001101110000;
		16'b0001110000001000 : data_out =  24'b000000100001001111111000;
		16'b0001110000001010 : data_out =  24'b000000100001010010000000;
		16'b0001110000001100 : data_out =  24'b000000100001010100001001;
		16'b0001110000001110 : data_out =  24'b000000100001010110010001;
		16'b0001110000010000 : data_out =  24'b000000100001011000011010;
		16'b0001110000010010 : data_out =  24'b000000100001011010100011;
		16'b0001110000010100 : data_out =  24'b000000100001011100101100;
		16'b0001110000010110 : data_out =  24'b000000100001011110110101;
		16'b0001110000011000 : data_out =  24'b000000100001100000111110;
		16'b0001110000011010 : data_out =  24'b000000100001100011000111;
		16'b0001110000011100 : data_out =  24'b000000100001100101010001;
		16'b0001110000011110 : data_out =  24'b000000100001100111011010;
		16'b0001110000100000 : data_out =  24'b000000100001101001100100;
		16'b0001110000100010 : data_out =  24'b000000100001101011101110;
		16'b0001110000100100 : data_out =  24'b000000100001101101111000;
		16'b0001110000100110 : data_out =  24'b000000100001110000000010;
		16'b0001110000101000 : data_out =  24'b000000100001110010001101;
		16'b0001110000101011 : data_out =  24'b000000100001110100010111;
		16'b0001110000101101 : data_out =  24'b000000100001110110100010;
		16'b0001110000101111 : data_out =  24'b000000100001111000101100;
		16'b0001110000110001 : data_out =  24'b000000100001111010110111;
		16'b0001110000110011 : data_out =  24'b000000100001111101000010;
		16'b0001110000110101 : data_out =  24'b000000100001111111001101;
		16'b0001110000110111 : data_out =  24'b000000100010000001011001;
		16'b0001110000111001 : data_out =  24'b000000100010000011100100;
		16'b0001110000111011 : data_out =  24'b000000100010000101110000;
		16'b0001110000111101 : data_out =  24'b000000100010000111111011;
		16'b0001110000111111 : data_out =  24'b000000100010001010000111;
		16'b0001110001000001 : data_out =  24'b000000100010001100010011;
		16'b0001110001000011 : data_out =  24'b000000100010001110011111;
		16'b0001110001000101 : data_out =  24'b000000100010010000101011;
		16'b0001110001000111 : data_out =  24'b000000100010010010111000;
		16'b0001110001001001 : data_out =  24'b000000100010010101000100;
		16'b0001110001001011 : data_out =  24'b000000100010010111010001;
		16'b0001110001001101 : data_out =  24'b000000100010011001011110;
		16'b0001110001001111 : data_out =  24'b000000100010011011101011;
		16'b0001110001010001 : data_out =  24'b000000100010011101111000;
		16'b0001110001010011 : data_out =  24'b000000100010100000000101;
		16'b0001110001010110 : data_out =  24'b000000100010100010010011;
		16'b0001110001011000 : data_out =  24'b000000100010100100100000;
		16'b0001110001011010 : data_out =  24'b000000100010100110101110;
		16'b0001110001011100 : data_out =  24'b000000100010101000111100;
		16'b0001110001011110 : data_out =  24'b000000100010101011001010;
		16'b0001110001100000 : data_out =  24'b000000100010101101011000;
		16'b0001110001100010 : data_out =  24'b000000100010101111100110;
		16'b0001110001100100 : data_out =  24'b000000100010110001110100;
		16'b0001110001100110 : data_out =  24'b000000100010110100000011;
		16'b0001110001101000 : data_out =  24'b000000100010110110010010;
		16'b0001110001101010 : data_out =  24'b000000100010111000100000;
		16'b0001110001101100 : data_out =  24'b000000100010111010101111;
		16'b0001110001101110 : data_out =  24'b000000100010111100111110;
		16'b0001110001110000 : data_out =  24'b000000100010111111001110;
		16'b0001110001110010 : data_out =  24'b000000100011000001011101;
		16'b0001110001110100 : data_out =  24'b000000100011000011101101;
		16'b0001110001110110 : data_out =  24'b000000100011000101111100;
		16'b0001110001111000 : data_out =  24'b000000100011001000001100;
		16'b0001110001111010 : data_out =  24'b000000100011001010011100;
		16'b0001110001111100 : data_out =  24'b000000100011001100101100;
		16'b0001110001111110 : data_out =  24'b000000100011001110111100;
		16'b0001110010000001 : data_out =  24'b000000100011010001001101;
		16'b0001110010000011 : data_out =  24'b000000100011010011011101;
		16'b0001110010000101 : data_out =  24'b000000100011010101101110;
		16'b0001110010000111 : data_out =  24'b000000100011010111111111;
		16'b0001110010001001 : data_out =  24'b000000100011011010010000;
		16'b0001110010001011 : data_out =  24'b000000100011011100100001;
		16'b0001110010001101 : data_out =  24'b000000100011011110110010;
		16'b0001110010001111 : data_out =  24'b000000100011100001000011;
		16'b0001110010010001 : data_out =  24'b000000100011100011010101;
		16'b0001110010010011 : data_out =  24'b000000100011100101100111;
		16'b0001110010010101 : data_out =  24'b000000100011100111111001;
		16'b0001110010010111 : data_out =  24'b000000100011101010001011;
		16'b0001110010011001 : data_out =  24'b000000100011101100011101;
		16'b0001110010011011 : data_out =  24'b000000100011101110101111;
		16'b0001110010011101 : data_out =  24'b000000100011110001000001;
		16'b0001110010011111 : data_out =  24'b000000100011110011010100;
		16'b0001110010100001 : data_out =  24'b000000100011110101100111;
		16'b0001110010100011 : data_out =  24'b000000100011110111111010;
		16'b0001110010100101 : data_out =  24'b000000100011111010001101;
		16'b0001110010100111 : data_out =  24'b000000100011111100100000;
		16'b0001110010101001 : data_out =  24'b000000100011111110110011;
		16'b0001110010101100 : data_out =  24'b000000100100000001000110;
		16'b0001110010101110 : data_out =  24'b000000100100000011011010;
		16'b0001110010110000 : data_out =  24'b000000100100000101101110;
		16'b0001110010110010 : data_out =  24'b000000100100001000000010;
		16'b0001110010110100 : data_out =  24'b000000100100001010010110;
		16'b0001110010110110 : data_out =  24'b000000100100001100101010;
		16'b0001110010111000 : data_out =  24'b000000100100001110111110;
		16'b0001110010111010 : data_out =  24'b000000100100010001010011;
		16'b0001110010111100 : data_out =  24'b000000100100010011100111;
		16'b0001110010111110 : data_out =  24'b000000100100010101111100;
		16'b0001110011000000 : data_out =  24'b000000100100011000010001;
		16'b0001110011000010 : data_out =  24'b000000100100011010100110;
		16'b0001110011000100 : data_out =  24'b000000100100011100111011;
		16'b0001110011000110 : data_out =  24'b000000100100011111010001;
		16'b0001110011001000 : data_out =  24'b000000100100100001100110;
		16'b0001110011001010 : data_out =  24'b000000100100100011111100;
		16'b0001110011001100 : data_out =  24'b000000100100100110010010;
		16'b0001110011001110 : data_out =  24'b000000100100101000101000;
		16'b0001110011010000 : data_out =  24'b000000100100101010111110;
		16'b0001110011010010 : data_out =  24'b000000100100101101010100;
		16'b0001110011010100 : data_out =  24'b000000100100101111101011;
		16'b0001110011010111 : data_out =  24'b000000100100110010000001;
		16'b0001110011011001 : data_out =  24'b000000100100110100011000;
		16'b0001110011011011 : data_out =  24'b000000100100110110101111;
		16'b0001110011011101 : data_out =  24'b000000100100111001000110;
		16'b0001110011011111 : data_out =  24'b000000100100111011011101;
		16'b0001110011100001 : data_out =  24'b000000100100111101110100;
		16'b0001110011100011 : data_out =  24'b000000100101000000001100;
		16'b0001110011100101 : data_out =  24'b000000100101000010100100;
		16'b0001110011100111 : data_out =  24'b000000100101000100111011;
		16'b0001110011101001 : data_out =  24'b000000100101000111010011;
		16'b0001110011101011 : data_out =  24'b000000100101001001101011;
		16'b0001110011101101 : data_out =  24'b000000100101001100000100;
		16'b0001110011101111 : data_out =  24'b000000100101001110011100;
		16'b0001110011110001 : data_out =  24'b000000100101010000110101;
		16'b0001110011110011 : data_out =  24'b000000100101010011001101;
		16'b0001110011110101 : data_out =  24'b000000100101010101100110;
		16'b0001110011110111 : data_out =  24'b000000100101010111111111;
		16'b0001110011111001 : data_out =  24'b000000100101011010011000;
		16'b0001110011111011 : data_out =  24'b000000100101011100110010;
		16'b0001110011111101 : data_out =  24'b000000100101011111001011;
		16'b0001110011111111 : data_out =  24'b000000100101100001100101;
		16'b0001110100000010 : data_out =  24'b000000100101100011111111;
		16'b0001110100000100 : data_out =  24'b000000100101100110011000;
		16'b0001110100000110 : data_out =  24'b000000100101101000110011;
		16'b0001110100001000 : data_out =  24'b000000100101101011001101;
		16'b0001110100001010 : data_out =  24'b000000100101101101100111;
		16'b0001110100001100 : data_out =  24'b000000100101110000000010;
		16'b0001110100001110 : data_out =  24'b000000100101110010011100;
		16'b0001110100010000 : data_out =  24'b000000100101110100110111;
		16'b0001110100010010 : data_out =  24'b000000100101110111010010;
		16'b0001110100010100 : data_out =  24'b000000100101111001101101;
		16'b0001110100010110 : data_out =  24'b000000100101111100001001;
		16'b0001110100011000 : data_out =  24'b000000100101111110100100;
		16'b0001110100011010 : data_out =  24'b000000100110000001000000;
		16'b0001110100011100 : data_out =  24'b000000100110000011011100;
		16'b0001110100011110 : data_out =  24'b000000100110000101111000;
		16'b0001110100100000 : data_out =  24'b000000100110001000010100;
		16'b0001110100100010 : data_out =  24'b000000100110001010110000;
		16'b0001110100100100 : data_out =  24'b000000100110001101001100;
		16'b0001110100100110 : data_out =  24'b000000100110001111101001;
		16'b0001110100101000 : data_out =  24'b000000100110010010000110;
		16'b0001110100101011 : data_out =  24'b000000100110010100100011;
		16'b0001110100101101 : data_out =  24'b000000100110010111000000;
		16'b0001110100101111 : data_out =  24'b000000100110011001011101;
		16'b0001110100110001 : data_out =  24'b000000100110011011111010;
		16'b0001110100110011 : data_out =  24'b000000100110011110011000;
		16'b0001110100110101 : data_out =  24'b000000100110100000110101;
		16'b0001110100110111 : data_out =  24'b000000100110100011010011;
		16'b0001110100111001 : data_out =  24'b000000100110100101110001;
		16'b0001110100111011 : data_out =  24'b000000100110101000001111;
		16'b0001110100111101 : data_out =  24'b000000100110101010101110;
		16'b0001110100111111 : data_out =  24'b000000100110101101001100;
		16'b0001110101000001 : data_out =  24'b000000100110101111101011;
		16'b0001110101000011 : data_out =  24'b000000100110110010001010;
		16'b0001110101000101 : data_out =  24'b000000100110110100101000;
		16'b0001110101000111 : data_out =  24'b000000100110110111001000;
		16'b0001110101001001 : data_out =  24'b000000100110111001100111;
		16'b0001110101001011 : data_out =  24'b000000100110111100000110;
		16'b0001110101001101 : data_out =  24'b000000100110111110100110;
		16'b0001110101001111 : data_out =  24'b000000100111000001000110;
		16'b0001110101010001 : data_out =  24'b000000100111000011100101;
		16'b0001110101010011 : data_out =  24'b000000100111000110000101;
		16'b0001110101010110 : data_out =  24'b000000100111001000100110;
		16'b0001110101011000 : data_out =  24'b000000100111001011000110;
		16'b0001110101011010 : data_out =  24'b000000100111001101100111;
		16'b0001110101011100 : data_out =  24'b000000100111010000000111;
		16'b0001110101011110 : data_out =  24'b000000100111010010101000;
		16'b0001110101100000 : data_out =  24'b000000100111010101001001;
		16'b0001110101100010 : data_out =  24'b000000100111010111101010;
		16'b0001110101100100 : data_out =  24'b000000100111011010001100;
		16'b0001110101100110 : data_out =  24'b000000100111011100101101;
		16'b0001110101101000 : data_out =  24'b000000100111011111001111;
		16'b0001110101101010 : data_out =  24'b000000100111100001110001;
		16'b0001110101101100 : data_out =  24'b000000100111100100010011;
		16'b0001110101101110 : data_out =  24'b000000100111100110110101;
		16'b0001110101110000 : data_out =  24'b000000100111101001010111;
		16'b0001110101110010 : data_out =  24'b000000100111101011111010;
		16'b0001110101110100 : data_out =  24'b000000100111101110011100;
		16'b0001110101110110 : data_out =  24'b000000100111110000111111;
		16'b0001110101111000 : data_out =  24'b000000100111110011100010;
		16'b0001110101111010 : data_out =  24'b000000100111110110000101;
		16'b0001110101111100 : data_out =  24'b000000100111111000101000;
		16'b0001110101111110 : data_out =  24'b000000100111111011001100;
		16'b0001110110000001 : data_out =  24'b000000100111111101101111;
		16'b0001110110000011 : data_out =  24'b000000101000000000010011;
		16'b0001110110000101 : data_out =  24'b000000101000000010110111;
		16'b0001110110000111 : data_out =  24'b000000101000000101011011;
		16'b0001110110001001 : data_out =  24'b000000101000001000000000;
		16'b0001110110001011 : data_out =  24'b000000101000001010100100;
		16'b0001110110001101 : data_out =  24'b000000101000001101001001;
		16'b0001110110001111 : data_out =  24'b000000101000001111101101;
		16'b0001110110010001 : data_out =  24'b000000101000010010010010;
		16'b0001110110010011 : data_out =  24'b000000101000010100110111;
		16'b0001110110010101 : data_out =  24'b000000101000010111011101;
		16'b0001110110010111 : data_out =  24'b000000101000011010000010;
		16'b0001110110011001 : data_out =  24'b000000101000011100101000;
		16'b0001110110011011 : data_out =  24'b000000101000011111001101;
		16'b0001110110011101 : data_out =  24'b000000101000100001110011;
		16'b0001110110011111 : data_out =  24'b000000101000100100011001;
		16'b0001110110100001 : data_out =  24'b000000101000100111000000;
		16'b0001110110100011 : data_out =  24'b000000101000101001100110;
		16'b0001110110100101 : data_out =  24'b000000101000101100001101;
		16'b0001110110100111 : data_out =  24'b000000101000101110110011;
		16'b0001110110101001 : data_out =  24'b000000101000110001011010;
		16'b0001110110101100 : data_out =  24'b000000101000110100000001;
		16'b0001110110101110 : data_out =  24'b000000101000110110101001;
		16'b0001110110110000 : data_out =  24'b000000101000111001010000;
		16'b0001110110110010 : data_out =  24'b000000101000111011111000;
		16'b0001110110110100 : data_out =  24'b000000101000111110011111;
		16'b0001110110110110 : data_out =  24'b000000101001000001000111;
		16'b0001110110111000 : data_out =  24'b000000101001000011101111;
		16'b0001110110111010 : data_out =  24'b000000101001000110011000;
		16'b0001110110111100 : data_out =  24'b000000101001001001000000;
		16'b0001110110111110 : data_out =  24'b000000101001001011101001;
		16'b0001110111000000 : data_out =  24'b000000101001001110010010;
		16'b0001110111000010 : data_out =  24'b000000101001010000111010;
		16'b0001110111000100 : data_out =  24'b000000101001010011100100;
		16'b0001110111000110 : data_out =  24'b000000101001010110001101;
		16'b0001110111001000 : data_out =  24'b000000101001011000110110;
		16'b0001110111001010 : data_out =  24'b000000101001011011100000;
		16'b0001110111001100 : data_out =  24'b000000101001011110001010;
		16'b0001110111001110 : data_out =  24'b000000101001100000110100;
		16'b0001110111010000 : data_out =  24'b000000101001100011011110;
		16'b0001110111010010 : data_out =  24'b000000101001100110001000;
		16'b0001110111010100 : data_out =  24'b000000101001101000110010;
		16'b0001110111010111 : data_out =  24'b000000101001101011011101;
		16'b0001110111011001 : data_out =  24'b000000101001101110001000;
		16'b0001110111011011 : data_out =  24'b000000101001110000110011;
		16'b0001110111011101 : data_out =  24'b000000101001110011011110;
		16'b0001110111011111 : data_out =  24'b000000101001110110001001;
		16'b0001110111100001 : data_out =  24'b000000101001111000110101;
		16'b0001110111100011 : data_out =  24'b000000101001111011100001;
		16'b0001110111100101 : data_out =  24'b000000101001111110001100;
		16'b0001110111100111 : data_out =  24'b000000101010000000111000;
		16'b0001110111101001 : data_out =  24'b000000101010000011100101;
		16'b0001110111101011 : data_out =  24'b000000101010000110010001;
		16'b0001110111101101 : data_out =  24'b000000101010001000111101;
		16'b0001110111101111 : data_out =  24'b000000101010001011101010;
		16'b0001110111110001 : data_out =  24'b000000101010001110010111;
		16'b0001110111110011 : data_out =  24'b000000101010010001000100;
		16'b0001110111110101 : data_out =  24'b000000101010010011110001;
		16'b0001110111110111 : data_out =  24'b000000101010010110011111;
		16'b0001110111111001 : data_out =  24'b000000101010011001001100;
		16'b0001110111111011 : data_out =  24'b000000101010011011111010;
		16'b0001110111111101 : data_out =  24'b000000101010011110101000;
		16'b0001110111111111 : data_out =  24'b000000101010100001010110;
		16'b0001111000000010 : data_out =  24'b000000101010100100000100;
		16'b0001111000000100 : data_out =  24'b000000101010100110110011;
		16'b0001111000000110 : data_out =  24'b000000101010101001100001;
		16'b0001111000001000 : data_out =  24'b000000101010101100010000;
		16'b0001111000001010 : data_out =  24'b000000101010101110111111;
		16'b0001111000001100 : data_out =  24'b000000101010110001101110;
		16'b0001111000001110 : data_out =  24'b000000101010110100011101;
		16'b0001111000010000 : data_out =  24'b000000101010110111001101;
		16'b0001111000010010 : data_out =  24'b000000101010111001111100;
		16'b0001111000010100 : data_out =  24'b000000101010111100101100;
		16'b0001111000010110 : data_out =  24'b000000101010111111011100;
		16'b0001111000011000 : data_out =  24'b000000101011000010001100;
		16'b0001111000011010 : data_out =  24'b000000101011000100111101;
		16'b0001111000011100 : data_out =  24'b000000101011000111101101;
		16'b0001111000011110 : data_out =  24'b000000101011001010011110;
		16'b0001111000100000 : data_out =  24'b000000101011001101001111;
		16'b0001111000100010 : data_out =  24'b000000101011010000000000;
		16'b0001111000100100 : data_out =  24'b000000101011010010110001;
		16'b0001111000100110 : data_out =  24'b000000101011010101100011;
		16'b0001111000101000 : data_out =  24'b000000101011011000010100;
		16'b0001111000101011 : data_out =  24'b000000101011011011000110;
		16'b0001111000101101 : data_out =  24'b000000101011011101111000;
		16'b0001111000101111 : data_out =  24'b000000101011100000101010;
		16'b0001111000110001 : data_out =  24'b000000101011100011011100;
		16'b0001111000110011 : data_out =  24'b000000101011100110001111;
		16'b0001111000110101 : data_out =  24'b000000101011101001000010;
		16'b0001111000110111 : data_out =  24'b000000101011101011110100;
		16'b0001111000111001 : data_out =  24'b000000101011101110100111;
		16'b0001111000111011 : data_out =  24'b000000101011110001011011;
		16'b0001111000111101 : data_out =  24'b000000101011110100001110;
		16'b0001111000111111 : data_out =  24'b000000101011110111000010;
		16'b0001111001000001 : data_out =  24'b000000101011111001110101;
		16'b0001111001000011 : data_out =  24'b000000101011111100101001;
		16'b0001111001000101 : data_out =  24'b000000101011111111011101;
		16'b0001111001000111 : data_out =  24'b000000101100000010010010;
		16'b0001111001001001 : data_out =  24'b000000101100000101000110;
		16'b0001111001001011 : data_out =  24'b000000101100000111111011;
		16'b0001111001001101 : data_out =  24'b000000101100001010110000;
		16'b0001111001001111 : data_out =  24'b000000101100001101100101;
		16'b0001111001010001 : data_out =  24'b000000101100010000011010;
		16'b0001111001010011 : data_out =  24'b000000101100010011001111;
		16'b0001111001010110 : data_out =  24'b000000101100010110000101;
		16'b0001111001011000 : data_out =  24'b000000101100011000111010;
		16'b0001111001011010 : data_out =  24'b000000101100011011110000;
		16'b0001111001011100 : data_out =  24'b000000101100011110100110;
		16'b0001111001011110 : data_out =  24'b000000101100100001011101;
		16'b0001111001100000 : data_out =  24'b000000101100100100010011;
		16'b0001111001100010 : data_out =  24'b000000101100100111001010;
		16'b0001111001100100 : data_out =  24'b000000101100101010000001;
		16'b0001111001100110 : data_out =  24'b000000101100101100111000;
		16'b0001111001101000 : data_out =  24'b000000101100101111101111;
		16'b0001111001101010 : data_out =  24'b000000101100110010100110;
		16'b0001111001101100 : data_out =  24'b000000101100110101011110;
		16'b0001111001101110 : data_out =  24'b000000101100111000010101;
		16'b0001111001110000 : data_out =  24'b000000101100111011001101;
		16'b0001111001110010 : data_out =  24'b000000101100111110000101;
		16'b0001111001110100 : data_out =  24'b000000101101000000111110;
		16'b0001111001110110 : data_out =  24'b000000101101000011110110;
		16'b0001111001111000 : data_out =  24'b000000101101000110101111;
		16'b0001111001111010 : data_out =  24'b000000101101001001101000;
		16'b0001111001111100 : data_out =  24'b000000101101001100100001;
		16'b0001111001111110 : data_out =  24'b000000101101001111011010;
		16'b0001111010000001 : data_out =  24'b000000101101010010010011;
		16'b0001111010000011 : data_out =  24'b000000101101010101001101;
		16'b0001111010000101 : data_out =  24'b000000101101011000000111;
		16'b0001111010000111 : data_out =  24'b000000101101011011000001;
		16'b0001111010001001 : data_out =  24'b000000101101011101111011;
		16'b0001111010001011 : data_out =  24'b000000101101100000110101;
		16'b0001111010001101 : data_out =  24'b000000101101100011110000;
		16'b0001111010001111 : data_out =  24'b000000101101100110101010;
		16'b0001111010010001 : data_out =  24'b000000101101101001100101;
		16'b0001111010010011 : data_out =  24'b000000101101101100100000;
		16'b0001111010010101 : data_out =  24'b000000101101101111011100;
		16'b0001111010010111 : data_out =  24'b000000101101110010010111;
		16'b0001111010011001 : data_out =  24'b000000101101110101010011;
		16'b0001111010011011 : data_out =  24'b000000101101111000001110;
		16'b0001111010011101 : data_out =  24'b000000101101111011001010;
		16'b0001111010011111 : data_out =  24'b000000101101111110000111;
		16'b0001111010100001 : data_out =  24'b000000101110000001000011;
		16'b0001111010100011 : data_out =  24'b000000101110000100000000;
		16'b0001111010100101 : data_out =  24'b000000101110000110111100;
		16'b0001111010100111 : data_out =  24'b000000101110001001111001;
		16'b0001111010101001 : data_out =  24'b000000101110001100110111;
		16'b0001111010101100 : data_out =  24'b000000101110001111110100;
		16'b0001111010101110 : data_out =  24'b000000101110010010110001;
		16'b0001111010110000 : data_out =  24'b000000101110010101101111;
		16'b0001111010110010 : data_out =  24'b000000101110011000101101;
		16'b0001111010110100 : data_out =  24'b000000101110011011101011;
		16'b0001111010110110 : data_out =  24'b000000101110011110101001;
		16'b0001111010111000 : data_out =  24'b000000101110100001101000;
		16'b0001111010111010 : data_out =  24'b000000101110100100100111;
		16'b0001111010111100 : data_out =  24'b000000101110100111100101;
		16'b0001111010111110 : data_out =  24'b000000101110101010100100;
		16'b0001111011000000 : data_out =  24'b000000101110101101100100;
		16'b0001111011000010 : data_out =  24'b000000101110110000100011;
		16'b0001111011000100 : data_out =  24'b000000101110110011100011;
		16'b0001111011000110 : data_out =  24'b000000101110110110100011;
		16'b0001111011001000 : data_out =  24'b000000101110111001100011;
		16'b0001111011001010 : data_out =  24'b000000101110111100100011;
		16'b0001111011001100 : data_out =  24'b000000101110111111100011;
		16'b0001111011001110 : data_out =  24'b000000101111000010100100;
		16'b0001111011010000 : data_out =  24'b000000101111000101100100;
		16'b0001111011010010 : data_out =  24'b000000101111001000100101;
		16'b0001111011010100 : data_out =  24'b000000101111001011100111;
		16'b0001111011010111 : data_out =  24'b000000101111001110101000;
		16'b0001111011011001 : data_out =  24'b000000101111010001101001;
		16'b0001111011011011 : data_out =  24'b000000101111010100101011;
		16'b0001111011011101 : data_out =  24'b000000101111010111101101;
		16'b0001111011011111 : data_out =  24'b000000101111011010101111;
		16'b0001111011100001 : data_out =  24'b000000101111011101110010;
		16'b0001111011100011 : data_out =  24'b000000101111100000110100;
		16'b0001111011100101 : data_out =  24'b000000101111100011110111;
		16'b0001111011100111 : data_out =  24'b000000101111100110111010;
		16'b0001111011101001 : data_out =  24'b000000101111101001111101;
		16'b0001111011101011 : data_out =  24'b000000101111101101000000;
		16'b0001111011101101 : data_out =  24'b000000101111110000000100;
		16'b0001111011101111 : data_out =  24'b000000101111110011000111;
		16'b0001111011110001 : data_out =  24'b000000101111110110001011;
		16'b0001111011110011 : data_out =  24'b000000101111111001001111;
		16'b0001111011110101 : data_out =  24'b000000101111111100010100;
		16'b0001111011110111 : data_out =  24'b000000101111111111011000;
		16'b0001111011111001 : data_out =  24'b000000110000000010011101;
		16'b0001111011111011 : data_out =  24'b000000110000000101100010;
		16'b0001111011111101 : data_out =  24'b000000110000001000100111;
		16'b0001111011111111 : data_out =  24'b000000110000001011101100;
		16'b0001111100000010 : data_out =  24'b000000110000001110110001;
		16'b0001111100000100 : data_out =  24'b000000110000010001110111;
		16'b0001111100000110 : data_out =  24'b000000110000010100111101;
		16'b0001111100001000 : data_out =  24'b000000110000011000000011;
		16'b0001111100001010 : data_out =  24'b000000110000011011001001;
		16'b0001111100001100 : data_out =  24'b000000110000011110010000;
		16'b0001111100001110 : data_out =  24'b000000110000100001010110;
		16'b0001111100010000 : data_out =  24'b000000110000100100011101;
		16'b0001111100010010 : data_out =  24'b000000110000100111100100;
		16'b0001111100010100 : data_out =  24'b000000110000101010101011;
		16'b0001111100010110 : data_out =  24'b000000110000101101110011;
		16'b0001111100011000 : data_out =  24'b000000110000110000111010;
		16'b0001111100011010 : data_out =  24'b000000110000110100000010;
		16'b0001111100011100 : data_out =  24'b000000110000110111001010;
		16'b0001111100011110 : data_out =  24'b000000110000111010010010;
		16'b0001111100100000 : data_out =  24'b000000110000111101011011;
		16'b0001111100100010 : data_out =  24'b000000110001000000100100;
		16'b0001111100100100 : data_out =  24'b000000110001000011101100;
		16'b0001111100100110 : data_out =  24'b000000110001000110110101;
		16'b0001111100101000 : data_out =  24'b000000110001001001111111;
		16'b0001111100101011 : data_out =  24'b000000110001001101001000;
		16'b0001111100101101 : data_out =  24'b000000110001010000010010;
		16'b0001111100101111 : data_out =  24'b000000110001010011011100;
		16'b0001111100110001 : data_out =  24'b000000110001010110100110;
		16'b0001111100110011 : data_out =  24'b000000110001011001110000;
		16'b0001111100110101 : data_out =  24'b000000110001011100111010;
		16'b0001111100110111 : data_out =  24'b000000110001100000000101;
		16'b0001111100111001 : data_out =  24'b000000110001100011010000;
		16'b0001111100111011 : data_out =  24'b000000110001100110011011;
		16'b0001111100111101 : data_out =  24'b000000110001101001100110;
		16'b0001111100111111 : data_out =  24'b000000110001101100110010;
		16'b0001111101000001 : data_out =  24'b000000110001101111111101;
		16'b0001111101000011 : data_out =  24'b000000110001110011001001;
		16'b0001111101000101 : data_out =  24'b000000110001110110010101;
		16'b0001111101000111 : data_out =  24'b000000110001111001100010;
		16'b0001111101001001 : data_out =  24'b000000110001111100101110;
		16'b0001111101001011 : data_out =  24'b000000110001111111111011;
		16'b0001111101001101 : data_out =  24'b000000110010000011001000;
		16'b0001111101001111 : data_out =  24'b000000110010000110010101;
		16'b0001111101010001 : data_out =  24'b000000110010001001100010;
		16'b0001111101010011 : data_out =  24'b000000110010001100110000;
		16'b0001111101010110 : data_out =  24'b000000110010001111111101;
		16'b0001111101011000 : data_out =  24'b000000110010010011001011;
		16'b0001111101011010 : data_out =  24'b000000110010010110011001;
		16'b0001111101011100 : data_out =  24'b000000110010011001101000;
		16'b0001111101011110 : data_out =  24'b000000110010011100110110;
		16'b0001111101100000 : data_out =  24'b000000110010100000000101;
		16'b0001111101100010 : data_out =  24'b000000110010100011010100;
		16'b0001111101100100 : data_out =  24'b000000110010100110100011;
		16'b0001111101100110 : data_out =  24'b000000110010101001110011;
		16'b0001111101101000 : data_out =  24'b000000110010101101000010;
		16'b0001111101101010 : data_out =  24'b000000110010110000010010;
		16'b0001111101101100 : data_out =  24'b000000110010110011100010;
		16'b0001111101101110 : data_out =  24'b000000110010110110110010;
		16'b0001111101110000 : data_out =  24'b000000110010111010000010;
		16'b0001111101110010 : data_out =  24'b000000110010111101010011;
		16'b0001111101110100 : data_out =  24'b000000110011000000100100;
		16'b0001111101110110 : data_out =  24'b000000110011000011110101;
		16'b0001111101111000 : data_out =  24'b000000110011000111000110;
		16'b0001111101111010 : data_out =  24'b000000110011001010011000;
		16'b0001111101111100 : data_out =  24'b000000110011001101101001;
		16'b0001111101111110 : data_out =  24'b000000110011010000111011;
		16'b0001111110000001 : data_out =  24'b000000110011010100001101;
		16'b0001111110000011 : data_out =  24'b000000110011010111100000;
		16'b0001111110000101 : data_out =  24'b000000110011011010110010;
		16'b0001111110000111 : data_out =  24'b000000110011011110000101;
		16'b0001111110001001 : data_out =  24'b000000110011100001011000;
		16'b0001111110001011 : data_out =  24'b000000110011100100101011;
		16'b0001111110001101 : data_out =  24'b000000110011100111111110;
		16'b0001111110001111 : data_out =  24'b000000110011101011010010;
		16'b0001111110010001 : data_out =  24'b000000110011101110100110;
		16'b0001111110010011 : data_out =  24'b000000110011110001111010;
		16'b0001111110010101 : data_out =  24'b000000110011110101001110;
		16'b0001111110010111 : data_out =  24'b000000110011111000100010;
		16'b0001111110011001 : data_out =  24'b000000110011111011110111;
		16'b0001111110011011 : data_out =  24'b000000110011111111001100;
		16'b0001111110011101 : data_out =  24'b000000110100000010100001;
		16'b0001111110011111 : data_out =  24'b000000110100000101110110;
		16'b0001111110100001 : data_out =  24'b000000110100001001001011;
		16'b0001111110100011 : data_out =  24'b000000110100001100100001;
		16'b0001111110100101 : data_out =  24'b000000110100001111110111;
		16'b0001111110100111 : data_out =  24'b000000110100010011001101;
		16'b0001111110101001 : data_out =  24'b000000110100010110100011;
		16'b0001111110101100 : data_out =  24'b000000110100011001111010;
		16'b0001111110101110 : data_out =  24'b000000110100011101010001;
		16'b0001111110110000 : data_out =  24'b000000110100100000101000;
		16'b0001111110110010 : data_out =  24'b000000110100100011111111;
		16'b0001111110110100 : data_out =  24'b000000110100100111010110;
		16'b0001111110110110 : data_out =  24'b000000110100101010101110;
		16'b0001111110111000 : data_out =  24'b000000110100101110000110;
		16'b0001111110111010 : data_out =  24'b000000110100110001011110;
		16'b0001111110111100 : data_out =  24'b000000110100110100110110;
		16'b0001111110111110 : data_out =  24'b000000110100111000001111;
		16'b0001111111000000 : data_out =  24'b000000110100111011100111;
		16'b0001111111000010 : data_out =  24'b000000110100111111000000;
		16'b0001111111000100 : data_out =  24'b000000110101000010011001;
		16'b0001111111000110 : data_out =  24'b000000110101000101110011;
		16'b0001111111001000 : data_out =  24'b000000110101001001001100;
		16'b0001111111001010 : data_out =  24'b000000110101001100100110;
		16'b0001111111001100 : data_out =  24'b000000110101010000000000;
		16'b0001111111001110 : data_out =  24'b000000110101010011011010;
		16'b0001111111010000 : data_out =  24'b000000110101010110110101;
		16'b0001111111010010 : data_out =  24'b000000110101011010001111;
		16'b0001111111010100 : data_out =  24'b000000110101011101101010;
		16'b0001111111010111 : data_out =  24'b000000110101100001000101;
		16'b0001111111011001 : data_out =  24'b000000110101100100100001;
		16'b0001111111011011 : data_out =  24'b000000110101100111111100;
		16'b0001111111011101 : data_out =  24'b000000110101101011011000;
		16'b0001111111011111 : data_out =  24'b000000110101101110110100;
		16'b0001111111100001 : data_out =  24'b000000110101110010010000;
		16'b0001111111100011 : data_out =  24'b000000110101110101101100;
		16'b0001111111100101 : data_out =  24'b000000110101111001001001;
		16'b0001111111100111 : data_out =  24'b000000110101111100100110;
		16'b0001111111101001 : data_out =  24'b000000110110000000000011;
		16'b0001111111101011 : data_out =  24'b000000110110000011100000;
		16'b0001111111101101 : data_out =  24'b000000110110000110111110;
		16'b0001111111101111 : data_out =  24'b000000110110001010011100;
		16'b0001111111110001 : data_out =  24'b000000110110001101111010;
		16'b0001111111110011 : data_out =  24'b000000110110010001011000;
		16'b0001111111110101 : data_out =  24'b000000110110010100110110;
		16'b0001111111110111 : data_out =  24'b000000110110011000010101;
		16'b0001111111111001 : data_out =  24'b000000110110011011110100;
		16'b0001111111111011 : data_out =  24'b000000110110011111010011;
		16'b0001111111111101 : data_out =  24'b000000110110100010110010;
		16'b0001111111111111 : data_out =  24'b000000110110100110010010;
		16'b0010000000000010 : data_out =  24'b000000110110101001110001;
		16'b0010000000000100 : data_out =  24'b000000110110101101010001;
		16'b0010000000000110 : data_out =  24'b000000110110110000110001;
		16'b0010000000001000 : data_out =  24'b000000110110110100010010;
		16'b0010000000001010 : data_out =  24'b000000110110110111110010;
		16'b0010000000001100 : data_out =  24'b000000110110111011010011;
		16'b0010000000001110 : data_out =  24'b000000110110111110110100;
		16'b0010000000010000 : data_out =  24'b000000110111000010010110;
		16'b0010000000010010 : data_out =  24'b000000110111000101110111;
		16'b0010000000010100 : data_out =  24'b000000110111001001011001;
		16'b0010000000010110 : data_out =  24'b000000110111001100111011;
		16'b0010000000011000 : data_out =  24'b000000110111010000011101;
		16'b0010000000011010 : data_out =  24'b000000110111010100000000;
		16'b0010000000011100 : data_out =  24'b000000110111010111100010;
		16'b0010000000011110 : data_out =  24'b000000110111011011000101;
		16'b0010000000100000 : data_out =  24'b000000110111011110101000;
		16'b0010000000100010 : data_out =  24'b000000110111100010001100;
		16'b0010000000100100 : data_out =  24'b000000110111100101101111;
		16'b0010000000100110 : data_out =  24'b000000110111101001010011;
		16'b0010000000101000 : data_out =  24'b000000110111101100110111;
		16'b0010000000101011 : data_out =  24'b000000110111110000011011;
		16'b0010000000101101 : data_out =  24'b000000110111110100000000;
		16'b0010000000101111 : data_out =  24'b000000110111110111100101;
		16'b0010000000110001 : data_out =  24'b000000110111111011001010;
		16'b0010000000110011 : data_out =  24'b000000110111111110101111;
		16'b0010000000110101 : data_out =  24'b000000111000000010010100;
		16'b0010000000110111 : data_out =  24'b000000111000000101111010;
		16'b0010000000111001 : data_out =  24'b000000111000001001100000;
		16'b0010000000111011 : data_out =  24'b000000111000001101000110;
		16'b0010000000111101 : data_out =  24'b000000111000010000101100;
		16'b0010000000111111 : data_out =  24'b000000111000010100010011;
		16'b0010000001000001 : data_out =  24'b000000111000010111111010;
		16'b0010000001000011 : data_out =  24'b000000111000011011100001;
		16'b0010000001000101 : data_out =  24'b000000111000011111001000;
		16'b0010000001000111 : data_out =  24'b000000111000100010101111;
		16'b0010000001001001 : data_out =  24'b000000111000100110010111;
		16'b0010000001001011 : data_out =  24'b000000111000101001111111;
		16'b0010000001001101 : data_out =  24'b000000111000101101100111;
		16'b0010000001001111 : data_out =  24'b000000111000110001010000;
		16'b0010000001010001 : data_out =  24'b000000111000110100111000;
		16'b0010000001010011 : data_out =  24'b000000111000111000100001;
		16'b0010000001010110 : data_out =  24'b000000111000111100001010;
		16'b0010000001011000 : data_out =  24'b000000111000111111110100;
		16'b0010000001011010 : data_out =  24'b000000111001000011011101;
		16'b0010000001011100 : data_out =  24'b000000111001000111000111;
		16'b0010000001011110 : data_out =  24'b000000111001001010110001;
		16'b0010000001100000 : data_out =  24'b000000111001001110011011;
		16'b0010000001100010 : data_out =  24'b000000111001010010000110;
		16'b0010000001100100 : data_out =  24'b000000111001010101110001;
		16'b0010000001100110 : data_out =  24'b000000111001011001011011;
		16'b0010000001101000 : data_out =  24'b000000111001011101000111;
		16'b0010000001101010 : data_out =  24'b000000111001100000110010;
		16'b0010000001101100 : data_out =  24'b000000111001100100011110;
		16'b0010000001101110 : data_out =  24'b000000111001101000001010;
		16'b0010000001110000 : data_out =  24'b000000111001101011110110;
		16'b0010000001110010 : data_out =  24'b000000111001101111100010;
		16'b0010000001110100 : data_out =  24'b000000111001110011001111;
		16'b0010000001110110 : data_out =  24'b000000111001110110111100;
		16'b0010000001111000 : data_out =  24'b000000111001111010101001;
		16'b0010000001111010 : data_out =  24'b000000111001111110010110;
		16'b0010000001111100 : data_out =  24'b000000111010000010000100;
		16'b0010000001111110 : data_out =  24'b000000111010000101110010;
		16'b0010000010000001 : data_out =  24'b000000111010001001100000;
		16'b0010000010000011 : data_out =  24'b000000111010001101001110;
		16'b0010000010000101 : data_out =  24'b000000111010010000111101;
		16'b0010000010000111 : data_out =  24'b000000111010010100101011;
		16'b0010000010001001 : data_out =  24'b000000111010011000011010;
		16'b0010000010001011 : data_out =  24'b000000111010011100001010;
		16'b0010000010001101 : data_out =  24'b000000111010011111111001;
		16'b0010000010001111 : data_out =  24'b000000111010100011101001;
		16'b0010000010010001 : data_out =  24'b000000111010100111011001;
		16'b0010000010010011 : data_out =  24'b000000111010101011001001;
		16'b0010000010010101 : data_out =  24'b000000111010101110111001;
		16'b0010000010010111 : data_out =  24'b000000111010110010101010;
		16'b0010000010011001 : data_out =  24'b000000111010110110011011;
		16'b0010000010011011 : data_out =  24'b000000111010111010001100;
		16'b0010000010011101 : data_out =  24'b000000111010111101111110;
		16'b0010000010011111 : data_out =  24'b000000111011000001101111;
		16'b0010000010100001 : data_out =  24'b000000111011000101100001;
		16'b0010000010100011 : data_out =  24'b000000111011001001010011;
		16'b0010000010100101 : data_out =  24'b000000111011001101000110;
		16'b0010000010100111 : data_out =  24'b000000111011010000111000;
		16'b0010000010101001 : data_out =  24'b000000111011010100101011;
		16'b0010000010101100 : data_out =  24'b000000111011011000011110;
		16'b0010000010101110 : data_out =  24'b000000111011011100010010;
		16'b0010000010110000 : data_out =  24'b000000111011100000000101;
		16'b0010000010110010 : data_out =  24'b000000111011100011111001;
		16'b0010000010110100 : data_out =  24'b000000111011100111101101;
		16'b0010000010110110 : data_out =  24'b000000111011101011100010;
		16'b0010000010111000 : data_out =  24'b000000111011101111010110;
		16'b0010000010111010 : data_out =  24'b000000111011110011001011;
		16'b0010000010111100 : data_out =  24'b000000111011110111000000;
		16'b0010000010111110 : data_out =  24'b000000111011111010110101;
		16'b0010000011000000 : data_out =  24'b000000111011111110101011;
		16'b0010000011000010 : data_out =  24'b000000111100000010100001;
		16'b0010000011000100 : data_out =  24'b000000111100000110010111;
		16'b0010000011000110 : data_out =  24'b000000111100001010001101;
		16'b0010000011001000 : data_out =  24'b000000111100001110000100;
		16'b0010000011001010 : data_out =  24'b000000111100010001111010;
		16'b0010000011001100 : data_out =  24'b000000111100010101110001;
		16'b0010000011001110 : data_out =  24'b000000111100011001101001;
		16'b0010000011010000 : data_out =  24'b000000111100011101100000;
		16'b0010000011010010 : data_out =  24'b000000111100100001011000;
		16'b0010000011010100 : data_out =  24'b000000111100100101010000;
		16'b0010000011010111 : data_out =  24'b000000111100101001001000;
		16'b0010000011011001 : data_out =  24'b000000111100101101000001;
		16'b0010000011011011 : data_out =  24'b000000111100110000111001;
		16'b0010000011011101 : data_out =  24'b000000111100110100110010;
		16'b0010000011011111 : data_out =  24'b000000111100111000101100;
		16'b0010000011100001 : data_out =  24'b000000111100111100100101;
		16'b0010000011100011 : data_out =  24'b000000111101000000011111;
		16'b0010000011100101 : data_out =  24'b000000111101000100011001;
		16'b0010000011100111 : data_out =  24'b000000111101001000010011;
		16'b0010000011101001 : data_out =  24'b000000111101001100001110;
		16'b0010000011101011 : data_out =  24'b000000111101010000001001;
		16'b0010000011101101 : data_out =  24'b000000111101010100000100;
		16'b0010000011101111 : data_out =  24'b000000111101010111111111;
		16'b0010000011110001 : data_out =  24'b000000111101011011111010;
		16'b0010000011110011 : data_out =  24'b000000111101011111110110;
		16'b0010000011110101 : data_out =  24'b000000111101100011110010;
		16'b0010000011110111 : data_out =  24'b000000111101100111101110;
		16'b0010000011111001 : data_out =  24'b000000111101101011101011;
		16'b0010000011111011 : data_out =  24'b000000111101101111101000;
		16'b0010000011111101 : data_out =  24'b000000111101110011100101;
		16'b0010000011111111 : data_out =  24'b000000111101110111100010;
		16'b0010000100000010 : data_out =  24'b000000111101111011100000;
		16'b0010000100000100 : data_out =  24'b000000111101111111011101;
		16'b0010000100000110 : data_out =  24'b000000111110000011011011;
		16'b0010000100001000 : data_out =  24'b000000111110000111011010;
		16'b0010000100001010 : data_out =  24'b000000111110001011011000;
		16'b0010000100001100 : data_out =  24'b000000111110001111010111;
		16'b0010000100001110 : data_out =  24'b000000111110010011010110;
		16'b0010000100010000 : data_out =  24'b000000111110010111010101;
		16'b0010000100010010 : data_out =  24'b000000111110011011010101;
		16'b0010000100010100 : data_out =  24'b000000111110011111010101;
		16'b0010000100010110 : data_out =  24'b000000111110100011010101;
		16'b0010000100011000 : data_out =  24'b000000111110100111010101;
		16'b0010000100011010 : data_out =  24'b000000111110101011010110;
		16'b0010000100011100 : data_out =  24'b000000111110101111010111;
		16'b0010000100011110 : data_out =  24'b000000111110110011011000;
		16'b0010000100100000 : data_out =  24'b000000111110110111011001;
		16'b0010000100100010 : data_out =  24'b000000111110111011011011;
		16'b0010000100100100 : data_out =  24'b000000111110111111011101;
		16'b0010000100100110 : data_out =  24'b000000111111000011011111;
		16'b0010000100101000 : data_out =  24'b000000111111000111100001;
		16'b0010000100101011 : data_out =  24'b000000111111001011100100;
		16'b0010000100101101 : data_out =  24'b000000111111001111100111;
		16'b0010000100101111 : data_out =  24'b000000111111010011101010;
		16'b0010000100110001 : data_out =  24'b000000111111010111101101;
		16'b0010000100110011 : data_out =  24'b000000111111011011110001;
		16'b0010000100110101 : data_out =  24'b000000111111011111110101;
		16'b0010000100110111 : data_out =  24'b000000111111100011111001;
		16'b0010000100111001 : data_out =  24'b000000111111100111111110;
		16'b0010000100111011 : data_out =  24'b000000111111101100000011;
		16'b0010000100111101 : data_out =  24'b000000111111110000001000;
		16'b0010000100111111 : data_out =  24'b000000111111110100001101;
		16'b0010000101000001 : data_out =  24'b000000111111111000010010;
		16'b0010000101000011 : data_out =  24'b000000111111111100011000;
		16'b0010000101000101 : data_out =  24'b000001000000000000011110;
		16'b0010000101000111 : data_out =  24'b000001000000000100100100;
		16'b0010000101001001 : data_out =  24'b000001000000001000101011;
		16'b0010000101001011 : data_out =  24'b000001000000001100110010;
		16'b0010000101001101 : data_out =  24'b000001000000010000111001;
		16'b0010000101001111 : data_out =  24'b000001000000010101000000;
		16'b0010000101010001 : data_out =  24'b000001000000011001001000;
		16'b0010000101010011 : data_out =  24'b000001000000011101010000;
		16'b0010000101010110 : data_out =  24'b000001000000100001011000;
		16'b0010000101011000 : data_out =  24'b000001000000100101100000;
		16'b0010000101011010 : data_out =  24'b000001000000101001101001;
		16'b0010000101011100 : data_out =  24'b000001000000101101110010;
		16'b0010000101011110 : data_out =  24'b000001000000110001111011;
		16'b0010000101100000 : data_out =  24'b000001000000110110000101;
		16'b0010000101100010 : data_out =  24'b000001000000111010001110;
		16'b0010000101100100 : data_out =  24'b000001000000111110011000;
		16'b0010000101100110 : data_out =  24'b000001000001000010100011;
		16'b0010000101101000 : data_out =  24'b000001000001000110101101;
		16'b0010000101101010 : data_out =  24'b000001000001001010111000;
		16'b0010000101101100 : data_out =  24'b000001000001001111000011;
		16'b0010000101101110 : data_out =  24'b000001000001010011001110;
		16'b0010000101110000 : data_out =  24'b000001000001010111011010;
		16'b0010000101110010 : data_out =  24'b000001000001011011100110;
		16'b0010000101110100 : data_out =  24'b000001000001011111110010;
		16'b0010000101110110 : data_out =  24'b000001000001100011111110;
		16'b0010000101111000 : data_out =  24'b000001000001101000001011;
		16'b0010000101111010 : data_out =  24'b000001000001101100011000;
		16'b0010000101111100 : data_out =  24'b000001000001110000100101;
		16'b0010000101111110 : data_out =  24'b000001000001110100110011;
		16'b0010000110000001 : data_out =  24'b000001000001111001000001;
		16'b0010000110000011 : data_out =  24'b000001000001111101001111;
		16'b0010000110000101 : data_out =  24'b000001000010000001011101;
		16'b0010000110000111 : data_out =  24'b000001000010000101101011;
		16'b0010000110001001 : data_out =  24'b000001000010001001111010;
		16'b0010000110001011 : data_out =  24'b000001000010001110001001;
		16'b0010000110001101 : data_out =  24'b000001000010010010011001;
		16'b0010000110001111 : data_out =  24'b000001000010010110101000;
		16'b0010000110010001 : data_out =  24'b000001000010011010111000;
		16'b0010000110010011 : data_out =  24'b000001000010011111001000;
		16'b0010000110010101 : data_out =  24'b000001000010100011011001;
		16'b0010000110010111 : data_out =  24'b000001000010100111101010;
		16'b0010000110011001 : data_out =  24'b000001000010101011111011;
		16'b0010000110011011 : data_out =  24'b000001000010110000001100;
		16'b0010000110011101 : data_out =  24'b000001000010110100011110;
		16'b0010000110011111 : data_out =  24'b000001000010111000101111;
		16'b0010000110100001 : data_out =  24'b000001000010111101000001;
		16'b0010000110100011 : data_out =  24'b000001000011000001010100;
		16'b0010000110100101 : data_out =  24'b000001000011000101100111;
		16'b0010000110100111 : data_out =  24'b000001000011001001111001;
		16'b0010000110101001 : data_out =  24'b000001000011001110001101;
		16'b0010000110101100 : data_out =  24'b000001000011010010100000;
		16'b0010000110101110 : data_out =  24'b000001000011010110110100;
		16'b0010000110110000 : data_out =  24'b000001000011011011001000;
		16'b0010000110110010 : data_out =  24'b000001000011011111011100;
		16'b0010000110110100 : data_out =  24'b000001000011100011110001;
		16'b0010000110110110 : data_out =  24'b000001000011101000000110;
		16'b0010000110111000 : data_out =  24'b000001000011101100011011;
		16'b0010000110111010 : data_out =  24'b000001000011110000110000;
		16'b0010000110111100 : data_out =  24'b000001000011110101000110;
		16'b0010000110111110 : data_out =  24'b000001000011111001011100;
		16'b0010000111000000 : data_out =  24'b000001000011111101110010;
		16'b0010000111000010 : data_out =  24'b000001000100000010001001;
		16'b0010000111000100 : data_out =  24'b000001000100000110011111;
		16'b0010000111000110 : data_out =  24'b000001000100001010110111;
		16'b0010000111001000 : data_out =  24'b000001000100001111001110;
		16'b0010000111001010 : data_out =  24'b000001000100010011100110;
		16'b0010000111001100 : data_out =  24'b000001000100010111111101;
		16'b0010000111001110 : data_out =  24'b000001000100011100010110;
		16'b0010000111010000 : data_out =  24'b000001000100100000101110;
		16'b0010000111010010 : data_out =  24'b000001000100100101000111;
		16'b0010000111010100 : data_out =  24'b000001000100101001100000;
		16'b0010000111010111 : data_out =  24'b000001000100101101111001;
		16'b0010000111011001 : data_out =  24'b000001000100110010010011;
		16'b0010000111011011 : data_out =  24'b000001000100110110101101;
		16'b0010000111011101 : data_out =  24'b000001000100111011000111;
		16'b0010000111011111 : data_out =  24'b000001000100111111100001;
		16'b0010000111100001 : data_out =  24'b000001000101000011111100;
		16'b0010000111100011 : data_out =  24'b000001000101001000010111;
		16'b0010000111100101 : data_out =  24'b000001000101001100110010;
		16'b0010000111100111 : data_out =  24'b000001000101010001001110;
		16'b0010000111101001 : data_out =  24'b000001000101010101101010;
		16'b0010000111101011 : data_out =  24'b000001000101011010000110;
		16'b0010000111101101 : data_out =  24'b000001000101011110100010;
		16'b0010000111101111 : data_out =  24'b000001000101100010111111;
		16'b0010000111110001 : data_out =  24'b000001000101100111011100;
		16'b0010000111110011 : data_out =  24'b000001000101101011111010;
		16'b0010000111110101 : data_out =  24'b000001000101110000010111;
		16'b0010000111110111 : data_out =  24'b000001000101110100110101;
		16'b0010000111111001 : data_out =  24'b000001000101111001010011;
		16'b0010000111111011 : data_out =  24'b000001000101111101110010;
		16'b0010000111111101 : data_out =  24'b000001000110000010010000;
		16'b0010000111111111 : data_out =  24'b000001000110000110101111;
		16'b0010001000000010 : data_out =  24'b000001000110001011001111;
		16'b0010001000000100 : data_out =  24'b000001000110001111101110;
		16'b0010001000000110 : data_out =  24'b000001000110010100001110;
		16'b0010001000001000 : data_out =  24'b000001000110011000101110;
		16'b0010001000001010 : data_out =  24'b000001000110011101001111;
		16'b0010001000001100 : data_out =  24'b000001000110100001101111;
		16'b0010001000001110 : data_out =  24'b000001000110100110010000;
		16'b0010001000010000 : data_out =  24'b000001000110101010110010;
		16'b0010001000010010 : data_out =  24'b000001000110101111010011;
		16'b0010001000010100 : data_out =  24'b000001000110110011110101;
		16'b0010001000010110 : data_out =  24'b000001000110111000010111;
		16'b0010001000011000 : data_out =  24'b000001000110111100111010;
		16'b0010001000011010 : data_out =  24'b000001000111000001011101;
		16'b0010001000011100 : data_out =  24'b000001000111000110000000;
		16'b0010001000011110 : data_out =  24'b000001000111001010100011;
		16'b0010001000100000 : data_out =  24'b000001000111001111000111;
		16'b0010001000100010 : data_out =  24'b000001000111010011101011;
		16'b0010001000100100 : data_out =  24'b000001000111011000001111;
		16'b0010001000100110 : data_out =  24'b000001000111011100110011;
		16'b0010001000101000 : data_out =  24'b000001000111100001011000;
		16'b0010001000101011 : data_out =  24'b000001000111100101111101;
		16'b0010001000101101 : data_out =  24'b000001000111101010100011;
		16'b0010001000101111 : data_out =  24'b000001000111101111001000;
		16'b0010001000110001 : data_out =  24'b000001000111110011101110;
		16'b0010001000110011 : data_out =  24'b000001000111111000010101;
		16'b0010001000110101 : data_out =  24'b000001000111111100111011;
		16'b0010001000110111 : data_out =  24'b000001001000000001100010;
		16'b0010001000111001 : data_out =  24'b000001001000000110001001;
		16'b0010001000111011 : data_out =  24'b000001001000001010110001;
		16'b0010001000111101 : data_out =  24'b000001001000001111011000;
		16'b0010001000111111 : data_out =  24'b000001001000010100000000;
		16'b0010001001000001 : data_out =  24'b000001001000011000101001;
		16'b0010001001000011 : data_out =  24'b000001001000011101010001;
		16'b0010001001000101 : data_out =  24'b000001001000100001111010;
		16'b0010001001000111 : data_out =  24'b000001001000100110100100;
		16'b0010001001001001 : data_out =  24'b000001001000101011001101;
		16'b0010001001001011 : data_out =  24'b000001001000101111110111;
		16'b0010001001001101 : data_out =  24'b000001001000110100100001;
		16'b0010001001001111 : data_out =  24'b000001001000111001001011;
		16'b0010001001010001 : data_out =  24'b000001001000111101110110;
		16'b0010001001010011 : data_out =  24'b000001001001000010100001;
		16'b0010001001010110 : data_out =  24'b000001001001000111001100;
		16'b0010001001011000 : data_out =  24'b000001001001001011111000;
		16'b0010001001011010 : data_out =  24'b000001001001010000100100;
		16'b0010001001011100 : data_out =  24'b000001001001010101010000;
		16'b0010001001011110 : data_out =  24'b000001001001011001111101;
		16'b0010001001100000 : data_out =  24'b000001001001011110101010;
		16'b0010001001100010 : data_out =  24'b000001001001100011010111;
		16'b0010001001100100 : data_out =  24'b000001001001101000000100;
		16'b0010001001100110 : data_out =  24'b000001001001101100110010;
		16'b0010001001101000 : data_out =  24'b000001001001110001100000;
		16'b0010001001101010 : data_out =  24'b000001001001110110001110;
		16'b0010001001101100 : data_out =  24'b000001001001111010111101;
		16'b0010001001101110 : data_out =  24'b000001001001111111101100;
		16'b0010001001110000 : data_out =  24'b000001001010000100011011;
		16'b0010001001110010 : data_out =  24'b000001001010001001001011;
		16'b0010001001110100 : data_out =  24'b000001001010001101111010;
		16'b0010001001110110 : data_out =  24'b000001001010010010101011;
		16'b0010001001111000 : data_out =  24'b000001001010010111011011;
		16'b0010001001111010 : data_out =  24'b000001001010011100001100;
		16'b0010001001111100 : data_out =  24'b000001001010100000111101;
		16'b0010001001111110 : data_out =  24'b000001001010100101101110;
		16'b0010001010000001 : data_out =  24'b000001001010101010100000;
		16'b0010001010000011 : data_out =  24'b000001001010101111010010;
		16'b0010001010000101 : data_out =  24'b000001001010110100000100;
		16'b0010001010000111 : data_out =  24'b000001001010111000110111;
		16'b0010001010001001 : data_out =  24'b000001001010111101101010;
		16'b0010001010001011 : data_out =  24'b000001001011000010011101;
		16'b0010001010001101 : data_out =  24'b000001001011000111010000;
		16'b0010001010001111 : data_out =  24'b000001001011001100000100;
		16'b0010001010010001 : data_out =  24'b000001001011010000111000;
		16'b0010001010010011 : data_out =  24'b000001001011010101101101;
		16'b0010001010010101 : data_out =  24'b000001001011011010100001;
		16'b0010001010010111 : data_out =  24'b000001001011011111010110;
		16'b0010001010011001 : data_out =  24'b000001001011100100001100;
		16'b0010001010011011 : data_out =  24'b000001001011101001000010;
		16'b0010001010011101 : data_out =  24'b000001001011101101110111;
		16'b0010001010011111 : data_out =  24'b000001001011110010101110;
		16'b0010001010100001 : data_out =  24'b000001001011110111100100;
		16'b0010001010100011 : data_out =  24'b000001001011111100011011;
		16'b0010001010100101 : data_out =  24'b000001001100000001010011;
		16'b0010001010100111 : data_out =  24'b000001001100000110001010;
		16'b0010001010101001 : data_out =  24'b000001001100001011000010;
		16'b0010001010101100 : data_out =  24'b000001001100001111111010;
		16'b0010001010101110 : data_out =  24'b000001001100010100110011;
		16'b0010001010110000 : data_out =  24'b000001001100011001101011;
		16'b0010001010110010 : data_out =  24'b000001001100011110100100;
		16'b0010001010110100 : data_out =  24'b000001001100100011011110;
		16'b0010001010110110 : data_out =  24'b000001001100101000011000;
		16'b0010001010111000 : data_out =  24'b000001001100101101010010;
		16'b0010001010111010 : data_out =  24'b000001001100110010001100;
		16'b0010001010111100 : data_out =  24'b000001001100110111000111;
		16'b0010001010111110 : data_out =  24'b000001001100111100000010;
		16'b0010001011000000 : data_out =  24'b000001001101000000111101;
		16'b0010001011000010 : data_out =  24'b000001001101000101111000;
		16'b0010001011000100 : data_out =  24'b000001001101001010110100;
		16'b0010001011000110 : data_out =  24'b000001001101001111110001;
		16'b0010001011001000 : data_out =  24'b000001001101010100101101;
		16'b0010001011001010 : data_out =  24'b000001001101011001101010;
		16'b0010001011001100 : data_out =  24'b000001001101011110100111;
		16'b0010001011001110 : data_out =  24'b000001001101100011100101;
		16'b0010001011010000 : data_out =  24'b000001001101101000100011;
		16'b0010001011010010 : data_out =  24'b000001001101101101100001;
		16'b0010001011010100 : data_out =  24'b000001001101110010011111;
		16'b0010001011010111 : data_out =  24'b000001001101110111011110;
		16'b0010001011011001 : data_out =  24'b000001001101111100011101;
		16'b0010001011011011 : data_out =  24'b000001001110000001011101;
		16'b0010001011011101 : data_out =  24'b000001001110000110011100;
		16'b0010001011011111 : data_out =  24'b000001001110001011011100;
		16'b0010001011100001 : data_out =  24'b000001001110010000011101;
		16'b0010001011100011 : data_out =  24'b000001001110010101011101;
		16'b0010001011100101 : data_out =  24'b000001001110011010011110;
		16'b0010001011100111 : data_out =  24'b000001001110011111100000;
		16'b0010001011101001 : data_out =  24'b000001001110100100100001;
		16'b0010001011101011 : data_out =  24'b000001001110101001100011;
		16'b0010001011101101 : data_out =  24'b000001001110101110100110;
		16'b0010001011101111 : data_out =  24'b000001001110110011101000;
		16'b0010001011110001 : data_out =  24'b000001001110111000101011;
		16'b0010001011110011 : data_out =  24'b000001001110111101101111;
		16'b0010001011110101 : data_out =  24'b000001001111000010110010;
		16'b0010001011110111 : data_out =  24'b000001001111000111110110;
		16'b0010001011111001 : data_out =  24'b000001001111001100111010;
		16'b0010001011111011 : data_out =  24'b000001001111010001111111;
		16'b0010001011111101 : data_out =  24'b000001001111010111000100;
		16'b0010001011111111 : data_out =  24'b000001001111011100001001;
		16'b0010001100000010 : data_out =  24'b000001001111100001001111;
		16'b0010001100000100 : data_out =  24'b000001001111100110010101;
		16'b0010001100000110 : data_out =  24'b000001001111101011011011;
		16'b0010001100001000 : data_out =  24'b000001001111110000100001;
		16'b0010001100001010 : data_out =  24'b000001001111110101101000;
		16'b0010001100001100 : data_out =  24'b000001001111111010101111;
		16'b0010001100001110 : data_out =  24'b000001001111111111110111;
		16'b0010001100010000 : data_out =  24'b000001010000000100111111;
		16'b0010001100010010 : data_out =  24'b000001010000001010000111;
		16'b0010001100010100 : data_out =  24'b000001010000001111001111;
		16'b0010001100010110 : data_out =  24'b000001010000010100011000;
		16'b0010001100011000 : data_out =  24'b000001010000011001100001;
		16'b0010001100011010 : data_out =  24'b000001010000011110101011;
		16'b0010001100011100 : data_out =  24'b000001010000100011110101;
		16'b0010001100011110 : data_out =  24'b000001010000101000111111;
		16'b0010001100100000 : data_out =  24'b000001010000101110001001;
		16'b0010001100100010 : data_out =  24'b000001010000110011010100;
		16'b0010001100100100 : data_out =  24'b000001010000111000011111;
		16'b0010001100100110 : data_out =  24'b000001010000111101101011;
		16'b0010001100101000 : data_out =  24'b000001010001000010110110;
		16'b0010001100101011 : data_out =  24'b000001010001001000000010;
		16'b0010001100101101 : data_out =  24'b000001010001001101001111;
		16'b0010001100101111 : data_out =  24'b000001010001010010011100;
		16'b0010001100110001 : data_out =  24'b000001010001010111101001;
		16'b0010001100110011 : data_out =  24'b000001010001011100110110;
		16'b0010001100110101 : data_out =  24'b000001010001100010000100;
		16'b0010001100110111 : data_out =  24'b000001010001100111010010;
		16'b0010001100111001 : data_out =  24'b000001010001101100100001;
		16'b0010001100111011 : data_out =  24'b000001010001110001101111;
		16'b0010001100111101 : data_out =  24'b000001010001110110111111;
		16'b0010001100111111 : data_out =  24'b000001010001111100001110;
		16'b0010001101000001 : data_out =  24'b000001010010000001011110;
		16'b0010001101000011 : data_out =  24'b000001010010000110101110;
		16'b0010001101000101 : data_out =  24'b000001010010001011111110;
		16'b0010001101000111 : data_out =  24'b000001010010010001001111;
		16'b0010001101001001 : data_out =  24'b000001010010010110100000;
		16'b0010001101001011 : data_out =  24'b000001010010011011110010;
		16'b0010001101001101 : data_out =  24'b000001010010100001000100;
		16'b0010001101001111 : data_out =  24'b000001010010100110010110;
		16'b0010001101010001 : data_out =  24'b000001010010101011101000;
		16'b0010001101010011 : data_out =  24'b000001010010110000111011;
		16'b0010001101010110 : data_out =  24'b000001010010110110001110;
		16'b0010001101011000 : data_out =  24'b000001010010111011100010;
		16'b0010001101011010 : data_out =  24'b000001010011000000110110;
		16'b0010001101011100 : data_out =  24'b000001010011000110001010;
		16'b0010001101011110 : data_out =  24'b000001010011001011011110;
		16'b0010001101100000 : data_out =  24'b000001010011010000110011;
		16'b0010001101100010 : data_out =  24'b000001010011010110001001;
		16'b0010001101100100 : data_out =  24'b000001010011011011011110;
		16'b0010001101100110 : data_out =  24'b000001010011100000110100;
		16'b0010001101101000 : data_out =  24'b000001010011100110001010;
		16'b0010001101101010 : data_out =  24'b000001010011101011100001;
		16'b0010001101101100 : data_out =  24'b000001010011110000111000;
		16'b0010001101101110 : data_out =  24'b000001010011110110001111;
		16'b0010001101110000 : data_out =  24'b000001010011111011100111;
		16'b0010001101110010 : data_out =  24'b000001010100000000111111;
		16'b0010001101110100 : data_out =  24'b000001010100000110010111;
		16'b0010001101110110 : data_out =  24'b000001010100001011101111;
		16'b0010001101111000 : data_out =  24'b000001010100010001001000;
		16'b0010001101111010 : data_out =  24'b000001010100010110100010;
		16'b0010001101111100 : data_out =  24'b000001010100011011111011;
		16'b0010001101111110 : data_out =  24'b000001010100100001010110;
		16'b0010001110000001 : data_out =  24'b000001010100100110110000;
		16'b0010001110000011 : data_out =  24'b000001010100101100001011;
		16'b0010001110000101 : data_out =  24'b000001010100110001100110;
		16'b0010001110000111 : data_out =  24'b000001010100110111000001;
		16'b0010001110001001 : data_out =  24'b000001010100111100011101;
		16'b0010001110001011 : data_out =  24'b000001010101000001111001;
		16'b0010001110001101 : data_out =  24'b000001010101000111010101;
		16'b0010001110001111 : data_out =  24'b000001010101001100110010;
		16'b0010001110010001 : data_out =  24'b000001010101010010001111;
		16'b0010001110010011 : data_out =  24'b000001010101010111101101;
		16'b0010001110010101 : data_out =  24'b000001010101011101001011;
		16'b0010001110010111 : data_out =  24'b000001010101100010101001;
		16'b0010001110011001 : data_out =  24'b000001010101101000000111;
		16'b0010001110011011 : data_out =  24'b000001010101101101100110;
		16'b0010001110011101 : data_out =  24'b000001010101110011000110;
		16'b0010001110011111 : data_out =  24'b000001010101111000100101;
		16'b0010001110100001 : data_out =  24'b000001010101111110000101;
		16'b0010001110100011 : data_out =  24'b000001010110000011100101;
		16'b0010001110100101 : data_out =  24'b000001010110001001000110;
		16'b0010001110100111 : data_out =  24'b000001010110001110100111;
		16'b0010001110101001 : data_out =  24'b000001010110010100001001;
		16'b0010001110101100 : data_out =  24'b000001010110011001101010;
		16'b0010001110101110 : data_out =  24'b000001010110011111001100;
		16'b0010001110110000 : data_out =  24'b000001010110100100101111;
		16'b0010001110110010 : data_out =  24'b000001010110101010010010;
		16'b0010001110110100 : data_out =  24'b000001010110101111110101;
		16'b0010001110110110 : data_out =  24'b000001010110110101011000;
		16'b0010001110111000 : data_out =  24'b000001010110111010111100;
		16'b0010001110111010 : data_out =  24'b000001010111000000100000;
		16'b0010001110111100 : data_out =  24'b000001010111000110000101;
		16'b0010001110111110 : data_out =  24'b000001010111001011101010;
		16'b0010001111000000 : data_out =  24'b000001010111010001001111;
		16'b0010001111000010 : data_out =  24'b000001010111010110110101;
		16'b0010001111000100 : data_out =  24'b000001010111011100011011;
		16'b0010001111000110 : data_out =  24'b000001010111100010000001;
		16'b0010001111001000 : data_out =  24'b000001010111100111101000;
		16'b0010001111001010 : data_out =  24'b000001010111101101001111;
		16'b0010001111001100 : data_out =  24'b000001010111110010110110;
		16'b0010001111001110 : data_out =  24'b000001010111111000011110;
		16'b0010001111010000 : data_out =  24'b000001010111111110000110;
		16'b0010001111010010 : data_out =  24'b000001011000000011101111;
		16'b0010001111010100 : data_out =  24'b000001011000001001010111;
		16'b0010001111010111 : data_out =  24'b000001011000001111000001;
		16'b0010001111011001 : data_out =  24'b000001011000010100101010;
		16'b0010001111011011 : data_out =  24'b000001011000011010010100;
		16'b0010001111011101 : data_out =  24'b000001011000011111111111;
		16'b0010001111011111 : data_out =  24'b000001011000100101101001;
		16'b0010001111100001 : data_out =  24'b000001011000101011010100;
		16'b0010001111100011 : data_out =  24'b000001011000110001000000;
		16'b0010001111100101 : data_out =  24'b000001011000110110101011;
		16'b0010001111100111 : data_out =  24'b000001011000111100011000;
		16'b0010001111101001 : data_out =  24'b000001011001000010000100;
		16'b0010001111101011 : data_out =  24'b000001011001000111110001;
		16'b0010001111101101 : data_out =  24'b000001011001001101011110;
		16'b0010001111101111 : data_out =  24'b000001011001010011001100;
		16'b0010001111110001 : data_out =  24'b000001011001011000111010;
		16'b0010001111110011 : data_out =  24'b000001011001011110101000;
		16'b0010001111110101 : data_out =  24'b000001011001100100010111;
		16'b0010001111110111 : data_out =  24'b000001011001101010000110;
		16'b0010001111111001 : data_out =  24'b000001011001101111110101;
		16'b0010001111111011 : data_out =  24'b000001011001110101100101;
		16'b0010001111111101 : data_out =  24'b000001011001111011010101;
		16'b0010001111111111 : data_out =  24'b000001011010000001000110;
		16'b0010010000000010 : data_out =  24'b000001011010000110110111;
		16'b0010010000000100 : data_out =  24'b000001011010001100101000;
		16'b0010010000000110 : data_out =  24'b000001011010010010011001;
		16'b0010010000001000 : data_out =  24'b000001011010011000001011;
		16'b0010010000001010 : data_out =  24'b000001011010011101111110;
		16'b0010010000001100 : data_out =  24'b000001011010100011110001;
		16'b0010010000001110 : data_out =  24'b000001011010101001100100;
		16'b0010010000010000 : data_out =  24'b000001011010101111010111;
		16'b0010010000010010 : data_out =  24'b000001011010110101001011;
		16'b0010010000010100 : data_out =  24'b000001011010111010111111;
		16'b0010010000010110 : data_out =  24'b000001011011000000110100;
		16'b0010010000011000 : data_out =  24'b000001011011000110101001;
		16'b0010010000011010 : data_out =  24'b000001011011001100011110;
		16'b0010010000011100 : data_out =  24'b000001011011010010010100;
		16'b0010010000011110 : data_out =  24'b000001011011011000001010;
		16'b0010010000100000 : data_out =  24'b000001011011011110000000;
		16'b0010010000100010 : data_out =  24'b000001011011100011110111;
		16'b0010010000100100 : data_out =  24'b000001011011101001101111;
		16'b0010010000100110 : data_out =  24'b000001011011101111100110;
		16'b0010010000101000 : data_out =  24'b000001011011110101011110;
		16'b0010010000101011 : data_out =  24'b000001011011111011010110;
		16'b0010010000101101 : data_out =  24'b000001011100000001001111;
		16'b0010010000101111 : data_out =  24'b000001011100000111001000;
		16'b0010010000110001 : data_out =  24'b000001011100001101000010;
		16'b0010010000110011 : data_out =  24'b000001011100010010111100;
		16'b0010010000110101 : data_out =  24'b000001011100011000110110;
		16'b0010010000110111 : data_out =  24'b000001011100011110110000;
		16'b0010010000111001 : data_out =  24'b000001011100100100101011;
		16'b0010010000111011 : data_out =  24'b000001011100101010100111;
		16'b0010010000111101 : data_out =  24'b000001011100110000100011;
		16'b0010010000111111 : data_out =  24'b000001011100110110011111;
		16'b0010010001000001 : data_out =  24'b000001011100111100011011;
		16'b0010010001000011 : data_out =  24'b000001011101000010011000;
		16'b0010010001000101 : data_out =  24'b000001011101001000010101;
		16'b0010010001000111 : data_out =  24'b000001011101001110010011;
		16'b0010010001001001 : data_out =  24'b000001011101010100010001;
		16'b0010010001001011 : data_out =  24'b000001011101011010001111;
		16'b0010010001001101 : data_out =  24'b000001011101100000001110;
		16'b0010010001001111 : data_out =  24'b000001011101100110001101;
		16'b0010010001010001 : data_out =  24'b000001011101101100001101;
		16'b0010010001010011 : data_out =  24'b000001011101110010001101;
		16'b0010010001010110 : data_out =  24'b000001011101111000001101;
		16'b0010010001011000 : data_out =  24'b000001011101111110001110;
		16'b0010010001011010 : data_out =  24'b000001011110000100001111;
		16'b0010010001011100 : data_out =  24'b000001011110001010010001;
		16'b0010010001011110 : data_out =  24'b000001011110010000010010;
		16'b0010010001100000 : data_out =  24'b000001011110010110010101;
		16'b0010010001100010 : data_out =  24'b000001011110011100010111;
		16'b0010010001100100 : data_out =  24'b000001011110100010011010;
		16'b0010010001100110 : data_out =  24'b000001011110101000011110;
		16'b0010010001101000 : data_out =  24'b000001011110101110100010;
		16'b0010010001101010 : data_out =  24'b000001011110110100100110;
		16'b0010010001101100 : data_out =  24'b000001011110111010101010;
		16'b0010010001101110 : data_out =  24'b000001011111000000101111;
		16'b0010010001110000 : data_out =  24'b000001011111000110110101;
		16'b0010010001110010 : data_out =  24'b000001011111001100111011;
		16'b0010010001110100 : data_out =  24'b000001011111010011000001;
		16'b0010010001110110 : data_out =  24'b000001011111011001000111;
		16'b0010010001111000 : data_out =  24'b000001011111011111001110;
		16'b0010010001111010 : data_out =  24'b000001011111100101010101;
		16'b0010010001111100 : data_out =  24'b000001011111101011011101;
		16'b0010010001111110 : data_out =  24'b000001011111110001100101;
		16'b0010010010000001 : data_out =  24'b000001011111110111101110;
		16'b0010010010000011 : data_out =  24'b000001011111111101110111;
		16'b0010010010000101 : data_out =  24'b000001100000000100000000;
		16'b0010010010000111 : data_out =  24'b000001100000001010001010;
		16'b0010010010001001 : data_out =  24'b000001100000010000010100;
		16'b0010010010001011 : data_out =  24'b000001100000010110011110;
		16'b0010010010001101 : data_out =  24'b000001100000011100101001;
		16'b0010010010001111 : data_out =  24'b000001100000100010110100;
		16'b0010010010010001 : data_out =  24'b000001100000101001000000;
		16'b0010010010010011 : data_out =  24'b000001100000101111001100;
		16'b0010010010010101 : data_out =  24'b000001100000110101011000;
		16'b0010010010010111 : data_out =  24'b000001100000111011100101;
		16'b0010010010011001 : data_out =  24'b000001100001000001110010;
		16'b0010010010011011 : data_out =  24'b000001100001001000000000;
		16'b0010010010011101 : data_out =  24'b000001100001001110001110;
		16'b0010010010011111 : data_out =  24'b000001100001010100011100;
		16'b0010010010100001 : data_out =  24'b000001100001011010101011;
		16'b0010010010100011 : data_out =  24'b000001100001100000111010;
		16'b0010010010100101 : data_out =  24'b000001100001100111001010;
		16'b0010010010100111 : data_out =  24'b000001100001101101011010;
		16'b0010010010101001 : data_out =  24'b000001100001110011101011;
		16'b0010010010101100 : data_out =  24'b000001100001111001111011;
		16'b0010010010101110 : data_out =  24'b000001100010000000001101;
		16'b0010010010110000 : data_out =  24'b000001100010000110011110;
		16'b0010010010110010 : data_out =  24'b000001100010001100110000;
		16'b0010010010110100 : data_out =  24'b000001100010010011000011;
		16'b0010010010110110 : data_out =  24'b000001100010011001010101;
		16'b0010010010111000 : data_out =  24'b000001100010011111101001;
		16'b0010010010111010 : data_out =  24'b000001100010100101111100;
		16'b0010010010111100 : data_out =  24'b000001100010101100010000;
		16'b0010010010111110 : data_out =  24'b000001100010110010100101;
		16'b0010010011000000 : data_out =  24'b000001100010111000111010;
		16'b0010010011000010 : data_out =  24'b000001100010111111001111;
		16'b0010010011000100 : data_out =  24'b000001100011000101100101;
		16'b0010010011000110 : data_out =  24'b000001100011001011111011;
		16'b0010010011001000 : data_out =  24'b000001100011010010010001;
		16'b0010010011001010 : data_out =  24'b000001100011011000101000;
		16'b0010010011001100 : data_out =  24'b000001100011011110111111;
		16'b0010010011001110 : data_out =  24'b000001100011100101010111;
		16'b0010010011010000 : data_out =  24'b000001100011101011101111;
		16'b0010010011010010 : data_out =  24'b000001100011110010001000;
		16'b0010010011010100 : data_out =  24'b000001100011111000100000;
		16'b0010010011010111 : data_out =  24'b000001100011111110111010;
		16'b0010010011011001 : data_out =  24'b000001100100000101010100;
		16'b0010010011011011 : data_out =  24'b000001100100001011101110;
		16'b0010010011011101 : data_out =  24'b000001100100010010001000;
		16'b0010010011011111 : data_out =  24'b000001100100011000100011;
		16'b0010010011100001 : data_out =  24'b000001100100011110111111;
		16'b0010010011100011 : data_out =  24'b000001100100100101011010;
		16'b0010010011100101 : data_out =  24'b000001100100101011110111;
		16'b0010010011100111 : data_out =  24'b000001100100110010010011;
		16'b0010010011101001 : data_out =  24'b000001100100111000110000;
		16'b0010010011101011 : data_out =  24'b000001100100111111001110;
		16'b0010010011101101 : data_out =  24'b000001100101000101101011;
		16'b0010010011101111 : data_out =  24'b000001100101001100001010;
		16'b0010010011110001 : data_out =  24'b000001100101010010101000;
		16'b0010010011110011 : data_out =  24'b000001100101011001001000;
		16'b0010010011110101 : data_out =  24'b000001100101011111100111;
		16'b0010010011110111 : data_out =  24'b000001100101100110000111;
		16'b0010010011111001 : data_out =  24'b000001100101101100100111;
		16'b0010010011111011 : data_out =  24'b000001100101110011001000;
		16'b0010010011111101 : data_out =  24'b000001100101111001101001;
		16'b0010010011111111 : data_out =  24'b000001100110000000001011;
		16'b0010010100000010 : data_out =  24'b000001100110000110101101;
		16'b0010010100000100 : data_out =  24'b000001100110001101001111;
		16'b0010010100000110 : data_out =  24'b000001100110010011110010;
		16'b0010010100001000 : data_out =  24'b000001100110011010010101;
		16'b0010010100001010 : data_out =  24'b000001100110100000111001;
		16'b0010010100001100 : data_out =  24'b000001100110100111011101;
		16'b0010010100001110 : data_out =  24'b000001100110101110000010;
		16'b0010010100010000 : data_out =  24'b000001100110110100100111;
		16'b0010010100010010 : data_out =  24'b000001100110111011001100;
		16'b0010010100010100 : data_out =  24'b000001100111000001110010;
		16'b0010010100010110 : data_out =  24'b000001100111001000011000;
		16'b0010010100011000 : data_out =  24'b000001100111001110111111;
		16'b0010010100011010 : data_out =  24'b000001100111010101100110;
		16'b0010010100011100 : data_out =  24'b000001100111011100001101;
		16'b0010010100011110 : data_out =  24'b000001100111100010110101;
		16'b0010010100100000 : data_out =  24'b000001100111101001011101;
		16'b0010010100100010 : data_out =  24'b000001100111110000000110;
		16'b0010010100100100 : data_out =  24'b000001100111110110101111;
		16'b0010010100100110 : data_out =  24'b000001100111111101011001;
		16'b0010010100101000 : data_out =  24'b000001101000000100000011;
		16'b0010010100101011 : data_out =  24'b000001101000001010101110;
		16'b0010010100101101 : data_out =  24'b000001101000010001011000;
		16'b0010010100101111 : data_out =  24'b000001101000011000000100;
		16'b0010010100110001 : data_out =  24'b000001101000011110101111;
		16'b0010010100110011 : data_out =  24'b000001101000100101011100;
		16'b0010010100110101 : data_out =  24'b000001101000101100001000;
		16'b0010010100110111 : data_out =  24'b000001101000110010110101;
		16'b0010010100111001 : data_out =  24'b000001101000111001100011;
		16'b0010010100111011 : data_out =  24'b000001101001000000010001;
		16'b0010010100111101 : data_out =  24'b000001101001000110111111;
		16'b0010010100111111 : data_out =  24'b000001101001001101101110;
		16'b0010010101000001 : data_out =  24'b000001101001010100011101;
		16'b0010010101000011 : data_out =  24'b000001101001011011001100;
		16'b0010010101000101 : data_out =  24'b000001101001100001111100;
		16'b0010010101000111 : data_out =  24'b000001101001101000101101;
		16'b0010010101001001 : data_out =  24'b000001101001101111011110;
		16'b0010010101001011 : data_out =  24'b000001101001110110001111;
		16'b0010010101001101 : data_out =  24'b000001101001111101000001;
		16'b0010010101001111 : data_out =  24'b000001101010000011110011;
		16'b0010010101010001 : data_out =  24'b000001101010001010100110;
		16'b0010010101010011 : data_out =  24'b000001101010010001011001;
		16'b0010010101010110 : data_out =  24'b000001101010011000001100;
		16'b0010010101011000 : data_out =  24'b000001101010011111000000;
		16'b0010010101011010 : data_out =  24'b000001101010100101110101;
		16'b0010010101011100 : data_out =  24'b000001101010101100101001;
		16'b0010010101011110 : data_out =  24'b000001101010110011011111;
		16'b0010010101100000 : data_out =  24'b000001101010111010010100;
		16'b0010010101100010 : data_out =  24'b000001101011000001001011;
		16'b0010010101100100 : data_out =  24'b000001101011001000000001;
		16'b0010010101100110 : data_out =  24'b000001101011001110111000;
		16'b0010010101101000 : data_out =  24'b000001101011010101110000;
		16'b0010010101101010 : data_out =  24'b000001101011011100100111;
		16'b0010010101101100 : data_out =  24'b000001101011100011100000;
		16'b0010010101101110 : data_out =  24'b000001101011101010011001;
		16'b0010010101110000 : data_out =  24'b000001101011110001010010;
		16'b0010010101110010 : data_out =  24'b000001101011111000001011;
		16'b0010010101110100 : data_out =  24'b000001101011111111000101;
		16'b0010010101110110 : data_out =  24'b000001101100000110000000;
		16'b0010010101111000 : data_out =  24'b000001101100001100111011;
		16'b0010010101111010 : data_out =  24'b000001101100010011110110;
		16'b0010010101111100 : data_out =  24'b000001101100011010110010;
		16'b0010010101111110 : data_out =  24'b000001101100100001101111;
		16'b0010010110000001 : data_out =  24'b000001101100101000101011;
		16'b0010010110000011 : data_out =  24'b000001101100101111101000;
		16'b0010010110000101 : data_out =  24'b000001101100110110100110;
		16'b0010010110000111 : data_out =  24'b000001101100111101100100;
		16'b0010010110001001 : data_out =  24'b000001101101000100100011;
		16'b0010010110001011 : data_out =  24'b000001101101001011100010;
		16'b0010010110001101 : data_out =  24'b000001101101010010100001;
		16'b0010010110001111 : data_out =  24'b000001101101011001100001;
		16'b0010010110010001 : data_out =  24'b000001101101100000100001;
		16'b0010010110010011 : data_out =  24'b000001101101100111100010;
		16'b0010010110010101 : data_out =  24'b000001101101101110100011;
		16'b0010010110010111 : data_out =  24'b000001101101110101100101;
		16'b0010010110011001 : data_out =  24'b000001101101111100100111;
		16'b0010010110011011 : data_out =  24'b000001101110000011101010;
		16'b0010010110011101 : data_out =  24'b000001101110001010101101;
		16'b0010010110011111 : data_out =  24'b000001101110010001110000;
		16'b0010010110100001 : data_out =  24'b000001101110011000110100;
		16'b0010010110100011 : data_out =  24'b000001101110011111111000;
		16'b0010010110100101 : data_out =  24'b000001101110100110111101;
		16'b0010010110100111 : data_out =  24'b000001101110101110000011;
		16'b0010010110101001 : data_out =  24'b000001101110110101001000;
		16'b0010010110101100 : data_out =  24'b000001101110111100001111;
		16'b0010010110101110 : data_out =  24'b000001101111000011010101;
		16'b0010010110110000 : data_out =  24'b000001101111001010011100;
		16'b0010010110110010 : data_out =  24'b000001101111010001100100;
		16'b0010010110110100 : data_out =  24'b000001101111011000101100;
		16'b0010010110110110 : data_out =  24'b000001101111011111110100;
		16'b0010010110111000 : data_out =  24'b000001101111100110111101;
		16'b0010010110111010 : data_out =  24'b000001101111101110000111;
		16'b0010010110111100 : data_out =  24'b000001101111110101010000;
		16'b0010010110111110 : data_out =  24'b000001101111111100011011;
		16'b0010010111000000 : data_out =  24'b000001110000000011100101;
		16'b0010010111000010 : data_out =  24'b000001110000001010110001;
		16'b0010010111000100 : data_out =  24'b000001110000010001111100;
		16'b0010010111000110 : data_out =  24'b000001110000011001001000;
		16'b0010010111001000 : data_out =  24'b000001110000100000010101;
		16'b0010010111001010 : data_out =  24'b000001110000100111100010;
		16'b0010010111001100 : data_out =  24'b000001110000101110110000;
		16'b0010010111001110 : data_out =  24'b000001110000110101111110;
		16'b0010010111010000 : data_out =  24'b000001110000111101001100;
		16'b0010010111010010 : data_out =  24'b000001110001000100011011;
		16'b0010010111010100 : data_out =  24'b000001110001001011101010;
		16'b0010010111010111 : data_out =  24'b000001110001010010111010;
		16'b0010010111011001 : data_out =  24'b000001110001011010001010;
		16'b0010010111011011 : data_out =  24'b000001110001100001011011;
		16'b0010010111011101 : data_out =  24'b000001110001101000101100;
		16'b0010010111011111 : data_out =  24'b000001110001101111111110;
		16'b0010010111100001 : data_out =  24'b000001110001110111010000;
		16'b0010010111100011 : data_out =  24'b000001110001111110100011;
		16'b0010010111100101 : data_out =  24'b000001110010000101110110;
		16'b0010010111100111 : data_out =  24'b000001110010001101001001;
		16'b0010010111101001 : data_out =  24'b000001110010010100011110;
		16'b0010010111101011 : data_out =  24'b000001110010011011110010;
		16'b0010010111101101 : data_out =  24'b000001110010100011000111;
		16'b0010010111101111 : data_out =  24'b000001110010101010011100;
		16'b0010010111110001 : data_out =  24'b000001110010110001110010;
		16'b0010010111110011 : data_out =  24'b000001110010111001001001;
		16'b0010010111110101 : data_out =  24'b000001110011000000011111;
		16'b0010010111110111 : data_out =  24'b000001110011000111110111;
		16'b0010010111111001 : data_out =  24'b000001110011001111001111;
		16'b0010010111111011 : data_out =  24'b000001110011010110100111;
		16'b0010010111111101 : data_out =  24'b000001110011011110000000;
		16'b0010010111111111 : data_out =  24'b000001110011100101011001;
		16'b0010011000000010 : data_out =  24'b000001110011101100110010;
		16'b0010011000000100 : data_out =  24'b000001110011110100001101;
		16'b0010011000000110 : data_out =  24'b000001110011111011100111;
		16'b0010011000001000 : data_out =  24'b000001110100000011000010;
		16'b0010011000001010 : data_out =  24'b000001110100001010011110;
		16'b0010011000001100 : data_out =  24'b000001110100010001111010;
		16'b0010011000001110 : data_out =  24'b000001110100011001010110;
		16'b0010011000010000 : data_out =  24'b000001110100100000110011;
		16'b0010011000010010 : data_out =  24'b000001110100101000010001;
		16'b0010011000010100 : data_out =  24'b000001110100101111101111;
		16'b0010011000010110 : data_out =  24'b000001110100110111001101;
		16'b0010011000011000 : data_out =  24'b000001110100111110101100;
		16'b0010011000011010 : data_out =  24'b000001110101000110001100;
		16'b0010011000011100 : data_out =  24'b000001110101001101101011;
		16'b0010011000011110 : data_out =  24'b000001110101010101001100;
		16'b0010011000100000 : data_out =  24'b000001110101011100101101;
		16'b0010011000100010 : data_out =  24'b000001110101100100001110;
		16'b0010011000100100 : data_out =  24'b000001110101101011110000;
		16'b0010011000100110 : data_out =  24'b000001110101110011010010;
		16'b0010011000101000 : data_out =  24'b000001110101111010110101;
		16'b0010011000101011 : data_out =  24'b000001110110000010011000;
		16'b0010011000101101 : data_out =  24'b000001110110001001111100;
		16'b0010011000101111 : data_out =  24'b000001110110010001100000;
		16'b0010011000110001 : data_out =  24'b000001110110011001000101;
		16'b0010011000110011 : data_out =  24'b000001110110100000101010;
		16'b0010011000110101 : data_out =  24'b000001110110101000001111;
		16'b0010011000110111 : data_out =  24'b000001110110101111110110;
		16'b0010011000111001 : data_out =  24'b000001110110110111011100;
		16'b0010011000111011 : data_out =  24'b000001110110111111000011;
		16'b0010011000111101 : data_out =  24'b000001110111000110101011;
		16'b0010011000111111 : data_out =  24'b000001110111001110010011;
		16'b0010011001000001 : data_out =  24'b000001110111010101111100;
		16'b0010011001000011 : data_out =  24'b000001110111011101100101;
		16'b0010011001000101 : data_out =  24'b000001110111100101001110;
		16'b0010011001000111 : data_out =  24'b000001110111101100111000;
		16'b0010011001001001 : data_out =  24'b000001110111110100100011;
		16'b0010011001001011 : data_out =  24'b000001110111111100001110;
		16'b0010011001001101 : data_out =  24'b000001111000000011111001;
		16'b0010011001001111 : data_out =  24'b000001111000001011100101;
		16'b0010011001010001 : data_out =  24'b000001111000010011010010;
		16'b0010011001010011 : data_out =  24'b000001111000011010111111;
		16'b0010011001010110 : data_out =  24'b000001111000100010101100;
		16'b0010011001011000 : data_out =  24'b000001111000101010011010;
		16'b0010011001011010 : data_out =  24'b000001111000110010001001;
		16'b0010011001011100 : data_out =  24'b000001111000111001111000;
		16'b0010011001011110 : data_out =  24'b000001111001000001100111;
		16'b0010011001100000 : data_out =  24'b000001111001001001010111;
		16'b0010011001100010 : data_out =  24'b000001111001010001001000;
		16'b0010011001100100 : data_out =  24'b000001111001011000111001;
		16'b0010011001100110 : data_out =  24'b000001111001100000101010;
		16'b0010011001101000 : data_out =  24'b000001111001101000011100;
		16'b0010011001101010 : data_out =  24'b000001111001110000001111;
		16'b0010011001101100 : data_out =  24'b000001111001111000000010;
		16'b0010011001101110 : data_out =  24'b000001111001111111110101;
		16'b0010011001110000 : data_out =  24'b000001111010000111101001;
		16'b0010011001110010 : data_out =  24'b000001111010001111011101;
		16'b0010011001110100 : data_out =  24'b000001111010010111010010;
		16'b0010011001110110 : data_out =  24'b000001111010011111001000;
		16'b0010011001111000 : data_out =  24'b000001111010100110111110;
		16'b0010011001111010 : data_out =  24'b000001111010101110110100;
		16'b0010011001111100 : data_out =  24'b000001111010110110101011;
		16'b0010011001111110 : data_out =  24'b000001111010111110100011;
		16'b0010011010000001 : data_out =  24'b000001111011000110011011;
		16'b0010011010000011 : data_out =  24'b000001111011001110010011;
		16'b0010011010000101 : data_out =  24'b000001111011010110001100;
		16'b0010011010000111 : data_out =  24'b000001111011011110000110;
		16'b0010011010001001 : data_out =  24'b000001111011100110000000;
		16'b0010011010001011 : data_out =  24'b000001111011101101111010;
		16'b0010011010001101 : data_out =  24'b000001111011110101110101;
		16'b0010011010001111 : data_out =  24'b000001111011111101110001;
		16'b0010011010010001 : data_out =  24'b000001111100000101101101;
		16'b0010011010010011 : data_out =  24'b000001111100001101101001;
		16'b0010011010010101 : data_out =  24'b000001111100010101100110;
		16'b0010011010010111 : data_out =  24'b000001111100011101100100;
		16'b0010011010011001 : data_out =  24'b000001111100100101100010;
		16'b0010011010011011 : data_out =  24'b000001111100101101100000;
		16'b0010011010011101 : data_out =  24'b000001111100110101011111;
		16'b0010011010011111 : data_out =  24'b000001111100111101011111;
		16'b0010011010100001 : data_out =  24'b000001111101000101011111;
		16'b0010011010100011 : data_out =  24'b000001111101001101100000;
		16'b0010011010100101 : data_out =  24'b000001111101010101100001;
		16'b0010011010100111 : data_out =  24'b000001111101011101100010;
		16'b0010011010101001 : data_out =  24'b000001111101100101100100;
		16'b0010011010101100 : data_out =  24'b000001111101101101100111;
		16'b0010011010101110 : data_out =  24'b000001111101110101101010;
		16'b0010011010110000 : data_out =  24'b000001111101111101101110;
		16'b0010011010110010 : data_out =  24'b000001111110000101110010;
		16'b0010011010110100 : data_out =  24'b000001111110001101110111;
		16'b0010011010110110 : data_out =  24'b000001111110010101111100;
		16'b0010011010111000 : data_out =  24'b000001111110011110000010;
		16'b0010011010111010 : data_out =  24'b000001111110100110001000;
		16'b0010011010111100 : data_out =  24'b000001111110101110001111;
		16'b0010011010111110 : data_out =  24'b000001111110110110010110;
		16'b0010011011000000 : data_out =  24'b000001111110111110011110;
		16'b0010011011000010 : data_out =  24'b000001111111000110100111;
		16'b0010011011000100 : data_out =  24'b000001111111001110101111;
		16'b0010011011000110 : data_out =  24'b000001111111010110111001;
		16'b0010011011001000 : data_out =  24'b000001111111011111000011;
		16'b0010011011001010 : data_out =  24'b000001111111100111001101;
		16'b0010011011001100 : data_out =  24'b000001111111101111011000;
		16'b0010011011001110 : data_out =  24'b000001111111110111100100;
		16'b0010011011010000 : data_out =  24'b000001111111111111110000;
		16'b0010011011010010 : data_out =  24'b000010000000000111111100;
		16'b0010011011010100 : data_out =  24'b000010000000010000001001;
		16'b0010011011010111 : data_out =  24'b000010000000011000010111;
		16'b0010011011011001 : data_out =  24'b000010000000100000100101;
		16'b0010011011011011 : data_out =  24'b000010000000101000110100;
		16'b0010011011011101 : data_out =  24'b000010000000110001000011;
		16'b0010011011011111 : data_out =  24'b000010000000111001010010;
		16'b0010011011100001 : data_out =  24'b000010000001000001100011;
		16'b0010011011100011 : data_out =  24'b000010000001001001110011;
		16'b0010011011100101 : data_out =  24'b000010000001010010000101;
		16'b0010011011100111 : data_out =  24'b000010000001011010010110;
		16'b0010011011101001 : data_out =  24'b000010000001100010101001;
		16'b0010011011101011 : data_out =  24'b000010000001101010111100;
		16'b0010011011101101 : data_out =  24'b000010000001110011001111;
		16'b0010011011101111 : data_out =  24'b000010000001111011100011;
		16'b0010011011110001 : data_out =  24'b000010000010000011110111;
		16'b0010011011110011 : data_out =  24'b000010000010001100001100;
		16'b0010011011110101 : data_out =  24'b000010000010010100100010;
		16'b0010011011110111 : data_out =  24'b000010000010011100111000;
		16'b0010011011111001 : data_out =  24'b000010000010100101001111;
		16'b0010011011111011 : data_out =  24'b000010000010101101100110;
		16'b0010011011111101 : data_out =  24'b000010000010110101111101;
		16'b0010011011111111 : data_out =  24'b000010000010111110010110;
		16'b0010011100000010 : data_out =  24'b000010000011000110101110;
		16'b0010011100000100 : data_out =  24'b000010000011001111001000;
		16'b0010011100000110 : data_out =  24'b000010000011010111100001;
		16'b0010011100001000 : data_out =  24'b000010000011011111111100;
		16'b0010011100001010 : data_out =  24'b000010000011101000010111;
		16'b0010011100001100 : data_out =  24'b000010000011110000110010;
		16'b0010011100001110 : data_out =  24'b000010000011111001001110;
		16'b0010011100010000 : data_out =  24'b000010000100000001101011;
		16'b0010011100010010 : data_out =  24'b000010000100001010001000;
		16'b0010011100010100 : data_out =  24'b000010000100010010100101;
		16'b0010011100010110 : data_out =  24'b000010000100011011000011;
		16'b0010011100011000 : data_out =  24'b000010000100100011100010;
		16'b0010011100011010 : data_out =  24'b000010000100101100000001;
		16'b0010011100011100 : data_out =  24'b000010000100110100100001;
		16'b0010011100011110 : data_out =  24'b000010000100111101000001;
		16'b0010011100100000 : data_out =  24'b000010000101000101100010;
		16'b0010011100100010 : data_out =  24'b000010000101001110000100;
		16'b0010011100100100 : data_out =  24'b000010000101010110100110;
		16'b0010011100100110 : data_out =  24'b000010000101011111001000;
		16'b0010011100101000 : data_out =  24'b000010000101100111101011;
		16'b0010011100101011 : data_out =  24'b000010000101110000001111;
		16'b0010011100101101 : data_out =  24'b000010000101111000110011;
		16'b0010011100101111 : data_out =  24'b000010000110000001010111;
		16'b0010011100110001 : data_out =  24'b000010000110001001111101;
		16'b0010011100110011 : data_out =  24'b000010000110010010100010;
		16'b0010011100110101 : data_out =  24'b000010000110011011001001;
		16'b0010011100110111 : data_out =  24'b000010000110100011110000;
		16'b0010011100111001 : data_out =  24'b000010000110101100010111;
		16'b0010011100111011 : data_out =  24'b000010000110110100111111;
		16'b0010011100111101 : data_out =  24'b000010000110111101101000;
		16'b0010011100111111 : data_out =  24'b000010000111000110010001;
		16'b0010011101000001 : data_out =  24'b000010000111001110111010;
		16'b0010011101000011 : data_out =  24'b000010000111010111100100;
		16'b0010011101000101 : data_out =  24'b000010000111100000001111;
		16'b0010011101000111 : data_out =  24'b000010000111101000111011;
		16'b0010011101001001 : data_out =  24'b000010000111110001100110;
		16'b0010011101001011 : data_out =  24'b000010000111111010010011;
		16'b0010011101001101 : data_out =  24'b000010001000000011000000;
		16'b0010011101001111 : data_out =  24'b000010001000001011101101;
		16'b0010011101010001 : data_out =  24'b000010001000010100011011;
		16'b0010011101010011 : data_out =  24'b000010001000011101001010;
		16'b0010011101010110 : data_out =  24'b000010001000100101111001;
		16'b0010011101011000 : data_out =  24'b000010001000101110101001;
		16'b0010011101011010 : data_out =  24'b000010001000110111011001;
		16'b0010011101011100 : data_out =  24'b000010001001000000001010;
		16'b0010011101011110 : data_out =  24'b000010001001001000111100;
		16'b0010011101100000 : data_out =  24'b000010001001010001101110;
		16'b0010011101100010 : data_out =  24'b000010001001011010100000;
		16'b0010011101100100 : data_out =  24'b000010001001100011010011;
		16'b0010011101100110 : data_out =  24'b000010001001101100000111;
		16'b0010011101101000 : data_out =  24'b000010001001110100111011;
		16'b0010011101101010 : data_out =  24'b000010001001111101110000;
		16'b0010011101101100 : data_out =  24'b000010001010000110100110;
		16'b0010011101101110 : data_out =  24'b000010001010001111011011;
		16'b0010011101110000 : data_out =  24'b000010001010011000010010;
		16'b0010011101110010 : data_out =  24'b000010001010100001001001;
		16'b0010011101110100 : data_out =  24'b000010001010101010000001;
		16'b0010011101110110 : data_out =  24'b000010001010110010111001;
		16'b0010011101111000 : data_out =  24'b000010001010111011110010;
		16'b0010011101111010 : data_out =  24'b000010001011000100101011;
		16'b0010011101111100 : data_out =  24'b000010001011001101100101;
		16'b0010011101111110 : data_out =  24'b000010001011010110100000;
		16'b0010011110000001 : data_out =  24'b000010001011011111011011;
		16'b0010011110000011 : data_out =  24'b000010001011101000010110;
		16'b0010011110000101 : data_out =  24'b000010001011110001010010;
		16'b0010011110000111 : data_out =  24'b000010001011111010001111;
		16'b0010011110001001 : data_out =  24'b000010001100000011001101;
		16'b0010011110001011 : data_out =  24'b000010001100001100001011;
		16'b0010011110001101 : data_out =  24'b000010001100010101001001;
		16'b0010011110001111 : data_out =  24'b000010001100011110001000;
		16'b0010011110010001 : data_out =  24'b000010001100100111001000;
		16'b0010011110010011 : data_out =  24'b000010001100110000001000;
		16'b0010011110010101 : data_out =  24'b000010001100111001001001;
		16'b0010011110010111 : data_out =  24'b000010001101000010001010;
		16'b0010011110011001 : data_out =  24'b000010001101001011001100;
		16'b0010011110011011 : data_out =  24'b000010001101010100001111;
		16'b0010011110011101 : data_out =  24'b000010001101011101010010;
		16'b0010011110011111 : data_out =  24'b000010001101100110010110;
		16'b0010011110100001 : data_out =  24'b000010001101101111011010;
		16'b0010011110100011 : data_out =  24'b000010001101111000011111;
		16'b0010011110100101 : data_out =  24'b000010001110000001100100;
		16'b0010011110100111 : data_out =  24'b000010001110001010101010;
		16'b0010011110101001 : data_out =  24'b000010001110010011110001;
		16'b0010011110101100 : data_out =  24'b000010001110011100111000;
		16'b0010011110101110 : data_out =  24'b000010001110100110000000;
		16'b0010011110110000 : data_out =  24'b000010001110101111001000;
		16'b0010011110110010 : data_out =  24'b000010001110111000010001;
		16'b0010011110110100 : data_out =  24'b000010001111000001011011;
		16'b0010011110110110 : data_out =  24'b000010001111001010100101;
		16'b0010011110111000 : data_out =  24'b000010001111010011101111;
		16'b0010011110111010 : data_out =  24'b000010001111011100111011;
		16'b0010011110111100 : data_out =  24'b000010001111100110000110;
		16'b0010011110111110 : data_out =  24'b000010001111101111010011;
		16'b0010011111000000 : data_out =  24'b000010001111111000100000;
		16'b0010011111000010 : data_out =  24'b000010010000000001101110;
		16'b0010011111000100 : data_out =  24'b000010010000001010111100;
		16'b0010011111000110 : data_out =  24'b000010010000010100001011;
		16'b0010011111001000 : data_out =  24'b000010010000011101011010;
		16'b0010011111001010 : data_out =  24'b000010010000100110101010;
		16'b0010011111001100 : data_out =  24'b000010010000101111111011;
		16'b0010011111001110 : data_out =  24'b000010010000111001001100;
		16'b0010011111010000 : data_out =  24'b000010010001000010011110;
		16'b0010011111010010 : data_out =  24'b000010010001001011110000;
		16'b0010011111010100 : data_out =  24'b000010010001010101000011;
		16'b0010011111010111 : data_out =  24'b000010010001011110010111;
		16'b0010011111011001 : data_out =  24'b000010010001100111101011;
		16'b0010011111011011 : data_out =  24'b000010010001110000111111;
		16'b0010011111011101 : data_out =  24'b000010010001111010010101;
		16'b0010011111011111 : data_out =  24'b000010010010000011101011;
		16'b0010011111100001 : data_out =  24'b000010010010001101000001;
		16'b0010011111100011 : data_out =  24'b000010010010010110011000;
		16'b0010011111100101 : data_out =  24'b000010010010011111110000;
		16'b0010011111100111 : data_out =  24'b000010010010101001001001;
		16'b0010011111101001 : data_out =  24'b000010010010110010100010;
		16'b0010011111101011 : data_out =  24'b000010010010111011111011;
		16'b0010011111101101 : data_out =  24'b000010010011000101010101;
		16'b0010011111101111 : data_out =  24'b000010010011001110110000;
		16'b0010011111110001 : data_out =  24'b000010010011011000001011;
		16'b0010011111110011 : data_out =  24'b000010010011100001100111;
		16'b0010011111110101 : data_out =  24'b000010010011101011000100;
		16'b0010011111110111 : data_out =  24'b000010010011110100100001;
		16'b0010011111111001 : data_out =  24'b000010010011111101111111;
		16'b0010011111111011 : data_out =  24'b000010010100000111011101;
		16'b0010011111111101 : data_out =  24'b000010010100010000111100;
	endcase
end
endmodule

